// Computer_System.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module Computer_System (
		inout  wire        av_config_SDAT,                                                          //                                                 av_config.SDAT
		output wire        av_config_SCLK,                                                          //                                                          .SCLK
		output wire        h2f_reset_reset_n,                                                       //                                                 h2f_reset.reset_n
		output wire        hps_io_hps_io_emac1_inst_TX_CLK,                                         //                                                    hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,                                           //                                                          .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,                                           //                                                          .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,                                           //                                                          .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,                                           //                                                          .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,                                           //                                                          .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,                                           //                                                          .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,                                            //                                                          .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL,                                         //                                                          .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL,                                         //                                                          .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK,                                         //                                                          .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,                                           //                                                          .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,                                           //                                                          .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,                                           //                                                          .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,                                             //                                                          .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,                                             //                                                          .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,                                             //                                                          .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,                                             //                                                          .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,                                             //                                                          .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,                                             //                                                          .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,                                             //                                                          .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,                                              //                                                          .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,                                              //                                                          .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,                                             //                                                          .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,                                              //                                                          .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,                                              //                                                          .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,                                              //                                                          .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,                                              //                                                          .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,                                              //                                                          .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,                                              //                                                          .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,                                              //                                                          .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,                                              //                                                          .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,                                              //                                                          .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,                                              //                                                          .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,                                             //                                                          .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,                                             //                                                          .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,                                             //                                                          .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,                                             //                                                          .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,                                            //                                                          .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,                                           //                                                          .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,                                           //                                                          .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,                                            //                                                          .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,                                             //                                                          .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,                                             //                                                          .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,                                             //                                                          .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,                                             //                                                          .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,                                             //                                                          .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,                                             //                                                          .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,                                          //                                                          .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,                                          //                                                          .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,                                          //                                                          .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO41,                                          //                                                          .hps_io_gpio_inst_GPIO41
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,                                          //                                                          .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,                                          //                                                          .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,                                          //                                                          .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,                                          //                                                          .hps_io_gpio_inst_GPIO61
		output wire [14:0] memory_mem_a,                                                            //                                                    memory.mem_a
		output wire [2:0]  memory_mem_ba,                                                           //                                                          .mem_ba
		output wire        memory_mem_ck,                                                           //                                                          .mem_ck
		output wire        memory_mem_ck_n,                                                         //                                                          .mem_ck_n
		output wire        memory_mem_cke,                                                          //                                                          .mem_cke
		output wire        memory_mem_cs_n,                                                         //                                                          .mem_cs_n
		output wire        memory_mem_ras_n,                                                        //                                                          .mem_ras_n
		output wire        memory_mem_cas_n,                                                        //                                                          .mem_cas_n
		output wire        memory_mem_we_n,                                                         //                                                          .mem_we_n
		output wire        memory_mem_reset_n,                                                      //                                                          .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                                                           //                                                          .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                                                          //                                                          .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                                                        //                                                          .mem_dqs_n
		output wire        memory_mem_odt,                                                          //                                                          .mem_odt
		output wire [3:0]  memory_mem_dm,                                                           //                                                          .mem_dm
		input  wire        memory_oct_rzqin,                                                        //                                                          .oct_rzqin
		output wire        pixel_clk_clk,                                                           //                                                 pixel_clk.clk
		output wire        pll_vga_clk_25_clk,                                                      //                                            pll_vga_clk_25.clk
		input  wire        rgba_image_sink_data_valid,                                              //                                           rgba_image_sink.data_valid
		input  wire [31:0] rgba_image_sink_input_data,                                              //                                                          .input_data
		input  wire [15:0] rgba_image_sink_img_width,                                               //                                                          .img_width
		input  wire [15:0] rgba_image_sink_img_height,                                              //                                                          .img_height
		output wire [31:0] rgba_image_src_data,                                                     //                                            rgba_image_src.data
		output wire        rgba_image_src_valid,                                                    //                                                          .valid
		input  wire        rgba_stream_reset_reset_n,                                               //                                         rgba_stream_reset.reset_n
		output wire [12:0] sdram_ctrl_addr,                                                         //                                                sdram_ctrl.addr
		output wire [1:0]  sdram_ctrl_ba,                                                           //                                                          .ba
		output wire        sdram_ctrl_cas_n,                                                        //                                                          .cas_n
		output wire        sdram_ctrl_cke,                                                          //                                                          .cke
		output wire        sdram_ctrl_cs_n,                                                         //                                                          .cs_n
		inout  wire [15:0] sdram_ctrl_dq,                                                           //                                                          .dq
		output wire [1:0]  sdram_ctrl_dqm,                                                          //                                                          .dqm
		output wire        sdram_ctrl_ras_n,                                                        //                                                          .ras_n
		output wire        sdram_ctrl_we_n,                                                         //                                                          .we_n
		input  wire        stream_control_endofpacket,                                              //                                            stream_control.endofpacket
		output wire        stream_control_ready,                                                    //                                                          .ready
		output wire        stream_control_sreset,                                                   //                                                          .sreset
		input  wire        system_pll_ref_clk_clk,                                                  //                                        system_pll_ref_clk.clk
		input  wire        system_pll_ref_reset_reset,                                              //                                      system_pll_ref_reset.reset
		input  wire        video_in_TD_CLK27,                                                       //                                                  video_in.TD_CLK27
		input  wire [7:0]  video_in_TD_DATA,                                                        //                                                          .TD_DATA
		input  wire        video_in_TD_HS,                                                          //                                                          .TD_HS
		input  wire        video_in_TD_VS,                                                          //                                                          .TD_VS
		input  wire        video_in_clk27_reset,                                                    //                                                          .clk27_reset
		output wire        video_in_TD_RESET,                                                       //                                                          .TD_RESET
		output wire        video_in_overflow_flag,                                                  //                                                          .overflow_flag
		input  wire [23:0] video_subsystem_video_in_feed_forward_avalon_forward_sink_data,          // video_subsystem_video_in_feed_forward_avalon_forward_sink.data
		input  wire        video_subsystem_video_in_feed_forward_avalon_forward_sink_startofpacket, //                                                          .startofpacket
		input  wire        video_subsystem_video_in_feed_forward_avalon_forward_sink_endofpacket,   //                                                          .endofpacket
		input  wire [1:0]  video_subsystem_video_in_feed_forward_avalon_forward_sink_empty,         //                                                          .empty
		input  wire        video_subsystem_video_in_feed_forward_avalon_forward_sink_valid,         //                                                          .valid
		output wire        video_subsystem_video_in_feed_forward_avalon_forward_sink_ready,         //                                                          .ready
		input  wire        video_subsystem_video_in_scaler_avalon_scaler_source_ready,              //      video_subsystem_video_in_scaler_avalon_scaler_source.ready
		output wire        video_subsystem_video_in_scaler_avalon_scaler_source_startofpacket,      //                                                          .startofpacket
		output wire        video_subsystem_video_in_scaler_avalon_scaler_source_endofpacket,        //                                                          .endofpacket
		output wire        video_subsystem_video_in_scaler_avalon_scaler_source_valid,              //                                                          .valid
		output wire [23:0] video_subsystem_video_in_scaler_avalon_scaler_source_data                //                                                          .data
	);

	wire          system_pll_reset_source_reset;                                  // System_PLL:reset_source_reset -> [PLL_VGA:rst, Video_Subsystem:reset_reset_n, rst_controller:reset_in0]
	wire          avalon_frame_writer_avalon_master_waitrequest;                  // mm_interconnect_0:Avalon_Frame_Writer_avalon_master_waitrequest -> Avalon_Frame_Writer:M_waitrequest
	wire   [31:0] avalon_frame_writer_avalon_master_address;                      // Avalon_Frame_Writer:M_address -> mm_interconnect_0:Avalon_Frame_Writer_avalon_master_address
	wire   [15:0] avalon_frame_writer_avalon_master_byteenable;                   // Avalon_Frame_Writer:M_byteenable -> mm_interconnect_0:Avalon_Frame_Writer_avalon_master_byteenable
	wire          avalon_frame_writer_avalon_master_write;                        // Avalon_Frame_Writer:M_write -> mm_interconnect_0:Avalon_Frame_Writer_avalon_master_write
	wire  [127:0] avalon_frame_writer_avalon_master_writedata;                    // Avalon_Frame_Writer:M_writedata -> mm_interconnect_0:Avalon_Frame_Writer_avalon_master_writedata
	wire    [6:0] avalon_frame_writer_avalon_master_burstcount;                   // Avalon_Frame_Writer:M_burstcount -> mm_interconnect_0:Avalon_Frame_Writer_avalon_master_burstcount
	wire          mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_waitrequest;       // ARM_A9_HPS:f2h_sdram1_WAITREQUEST -> mm_interconnect_0:ARM_A9_HPS_f2h_sdram1_data_waitrequest
	wire   [27:0] mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_address;           // mm_interconnect_0:ARM_A9_HPS_f2h_sdram1_data_address -> ARM_A9_HPS:f2h_sdram1_ADDRESS
	wire   [15:0] mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_byteenable;        // mm_interconnect_0:ARM_A9_HPS_f2h_sdram1_data_byteenable -> ARM_A9_HPS:f2h_sdram1_BYTEENABLE
	wire          mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_write;             // mm_interconnect_0:ARM_A9_HPS_f2h_sdram1_data_write -> ARM_A9_HPS:f2h_sdram1_WRITE
	wire  [127:0] mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_writedata;         // mm_interconnect_0:ARM_A9_HPS_f2h_sdram1_data_writedata -> ARM_A9_HPS:f2h_sdram1_WRITEDATA
	wire    [7:0] mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_burstcount;        // mm_interconnect_0:ARM_A9_HPS_f2h_sdram1_data_burstcount -> ARM_A9_HPS:f2h_sdram1_BURSTCOUNT
	wire          dot_product_avalon_master_waitrequest;                          // mm_interconnect_1:Dot_Product_avalon_master_waitrequest -> Dot_Product:master_waitrequest
	wire   [31:0] dot_product_avalon_master_readdata;                             // mm_interconnect_1:Dot_Product_avalon_master_readdata -> Dot_Product:master_readdata
	wire   [31:0] dot_product_avalon_master_address;                              // Dot_Product:master_address -> mm_interconnect_1:Dot_Product_avalon_master_address
	wire          dot_product_avalon_master_read;                                 // Dot_Product:master_read -> mm_interconnect_1:Dot_Product_avalon_master_read
	wire          dot_product_avalon_master_readdatavalid;                        // mm_interconnect_1:Dot_Product_avalon_master_readdatavalid -> Dot_Product:master_readdatavalid
	wire          dot_product_avalon_master_write;                                // Dot_Product:master_write -> mm_interconnect_1:Dot_Product_avalon_master_write
	wire   [31:0] dot_product_avalon_master_writedata;                            // Dot_Product:master_writedata -> mm_interconnect_1:Dot_Product_avalon_master_writedata
	wire    [1:0] arm_a9_hps_h2f_axi_master_awburst;                              // ARM_A9_HPS:h2f_AWBURST -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awburst
	wire    [3:0] arm_a9_hps_h2f_axi_master_arlen;                                // ARM_A9_HPS:h2f_ARLEN -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arlen
	wire   [15:0] arm_a9_hps_h2f_axi_master_wstrb;                                // ARM_A9_HPS:h2f_WSTRB -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_wstrb
	wire          arm_a9_hps_h2f_axi_master_wready;                               // mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_wready -> ARM_A9_HPS:h2f_WREADY
	wire   [11:0] arm_a9_hps_h2f_axi_master_rid;                                  // mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_rid -> ARM_A9_HPS:h2f_RID
	wire          arm_a9_hps_h2f_axi_master_rready;                               // ARM_A9_HPS:h2f_RREADY -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_rready
	wire    [3:0] arm_a9_hps_h2f_axi_master_awlen;                                // ARM_A9_HPS:h2f_AWLEN -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awlen
	wire   [11:0] arm_a9_hps_h2f_axi_master_wid;                                  // ARM_A9_HPS:h2f_WID -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_wid
	wire    [3:0] arm_a9_hps_h2f_axi_master_arcache;                              // ARM_A9_HPS:h2f_ARCACHE -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arcache
	wire          arm_a9_hps_h2f_axi_master_wvalid;                               // ARM_A9_HPS:h2f_WVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_wvalid
	wire   [29:0] arm_a9_hps_h2f_axi_master_araddr;                               // ARM_A9_HPS:h2f_ARADDR -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_araddr
	wire    [2:0] arm_a9_hps_h2f_axi_master_arprot;                               // ARM_A9_HPS:h2f_ARPROT -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arprot
	wire    [2:0] arm_a9_hps_h2f_axi_master_awprot;                               // ARM_A9_HPS:h2f_AWPROT -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awprot
	wire  [127:0] arm_a9_hps_h2f_axi_master_wdata;                                // ARM_A9_HPS:h2f_WDATA -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_wdata
	wire          arm_a9_hps_h2f_axi_master_arvalid;                              // ARM_A9_HPS:h2f_ARVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arvalid
	wire    [3:0] arm_a9_hps_h2f_axi_master_awcache;                              // ARM_A9_HPS:h2f_AWCACHE -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awcache
	wire   [11:0] arm_a9_hps_h2f_axi_master_arid;                                 // ARM_A9_HPS:h2f_ARID -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arid
	wire    [1:0] arm_a9_hps_h2f_axi_master_arlock;                               // ARM_A9_HPS:h2f_ARLOCK -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arlock
	wire    [1:0] arm_a9_hps_h2f_axi_master_awlock;                               // ARM_A9_HPS:h2f_AWLOCK -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awlock
	wire   [29:0] arm_a9_hps_h2f_axi_master_awaddr;                               // ARM_A9_HPS:h2f_AWADDR -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awaddr
	wire    [1:0] arm_a9_hps_h2f_axi_master_bresp;                                // mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_bresp -> ARM_A9_HPS:h2f_BRESP
	wire          arm_a9_hps_h2f_axi_master_arready;                              // mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arready -> ARM_A9_HPS:h2f_ARREADY
	wire  [127:0] arm_a9_hps_h2f_axi_master_rdata;                                // mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_rdata -> ARM_A9_HPS:h2f_RDATA
	wire          arm_a9_hps_h2f_axi_master_awready;                              // mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awready -> ARM_A9_HPS:h2f_AWREADY
	wire    [1:0] arm_a9_hps_h2f_axi_master_arburst;                              // ARM_A9_HPS:h2f_ARBURST -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arburst
	wire    [2:0] arm_a9_hps_h2f_axi_master_arsize;                               // ARM_A9_HPS:h2f_ARSIZE -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arsize
	wire          arm_a9_hps_h2f_axi_master_bready;                               // ARM_A9_HPS:h2f_BREADY -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_bready
	wire          arm_a9_hps_h2f_axi_master_rlast;                                // mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_rlast -> ARM_A9_HPS:h2f_RLAST
	wire          arm_a9_hps_h2f_axi_master_wlast;                                // ARM_A9_HPS:h2f_WLAST -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_wlast
	wire    [1:0] arm_a9_hps_h2f_axi_master_rresp;                                // mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_rresp -> ARM_A9_HPS:h2f_RRESP
	wire   [11:0] arm_a9_hps_h2f_axi_master_awid;                                 // ARM_A9_HPS:h2f_AWID -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awid
	wire   [11:0] arm_a9_hps_h2f_axi_master_bid;                                  // mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_bid -> ARM_A9_HPS:h2f_BID
	wire          arm_a9_hps_h2f_axi_master_bvalid;                               // mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_bvalid -> ARM_A9_HPS:h2f_BVALID
	wire    [2:0] arm_a9_hps_h2f_axi_master_awsize;                               // ARM_A9_HPS:h2f_AWSIZE -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awsize
	wire          arm_a9_hps_h2f_axi_master_awvalid;                              // ARM_A9_HPS:h2f_AWVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awvalid
	wire          arm_a9_hps_h2f_axi_master_rvalid;                               // mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_rvalid -> ARM_A9_HPS:h2f_RVALID
	wire          mm_interconnect_1_sram1_s1_chipselect;                          // mm_interconnect_1:SRAM1_s1_chipselect -> SRAM1:chipselect
	wire   [31:0] mm_interconnect_1_sram1_s1_readdata;                            // SRAM1:readdata -> mm_interconnect_1:SRAM1_s1_readdata
	wire    [9:0] mm_interconnect_1_sram1_s1_address;                             // mm_interconnect_1:SRAM1_s1_address -> SRAM1:address
	wire    [3:0] mm_interconnect_1_sram1_s1_byteenable;                          // mm_interconnect_1:SRAM1_s1_byteenable -> SRAM1:byteenable
	wire          mm_interconnect_1_sram1_s1_write;                               // mm_interconnect_1:SRAM1_s1_write -> SRAM1:write
	wire   [31:0] mm_interconnect_1_sram1_s1_writedata;                           // mm_interconnect_1:SRAM1_s1_writedata -> SRAM1:writedata
	wire          mm_interconnect_1_sram1_s1_clken;                               // mm_interconnect_1:SRAM1_s1_clken -> SRAM1:clken
	wire          mm_interconnect_1_sram2_s1_chipselect;                          // mm_interconnect_1:SRAM2_s1_chipselect -> SRAM2:chipselect
	wire   [31:0] mm_interconnect_1_sram2_s1_readdata;                            // SRAM2:readdata -> mm_interconnect_1:SRAM2_s1_readdata
	wire    [9:0] mm_interconnect_1_sram2_s1_address;                             // mm_interconnect_1:SRAM2_s1_address -> SRAM2:address
	wire    [3:0] mm_interconnect_1_sram2_s1_byteenable;                          // mm_interconnect_1:SRAM2_s1_byteenable -> SRAM2:byteenable
	wire          mm_interconnect_1_sram2_s1_write;                               // mm_interconnect_1:SRAM2_s1_write -> SRAM2:write
	wire   [31:0] mm_interconnect_1_sram2_s1_writedata;                           // mm_interconnect_1:SRAM2_s1_writedata -> SRAM2:writedata
	wire          mm_interconnect_1_sram2_s1_clken;                               // mm_interconnect_1:SRAM2_s1_clken -> SRAM2:clken
	wire          mm_interconnect_1_sdram_controller_s1_chipselect;               // mm_interconnect_1:SDRAM_Controller_s1_chipselect -> SDRAM_Controller:az_cs
	wire   [15:0] mm_interconnect_1_sdram_controller_s1_readdata;                 // SDRAM_Controller:za_data -> mm_interconnect_1:SDRAM_Controller_s1_readdata
	wire          mm_interconnect_1_sdram_controller_s1_waitrequest;              // SDRAM_Controller:za_waitrequest -> mm_interconnect_1:SDRAM_Controller_s1_waitrequest
	wire   [24:0] mm_interconnect_1_sdram_controller_s1_address;                  // mm_interconnect_1:SDRAM_Controller_s1_address -> SDRAM_Controller:az_addr
	wire          mm_interconnect_1_sdram_controller_s1_read;                     // mm_interconnect_1:SDRAM_Controller_s1_read -> SDRAM_Controller:az_rd_n
	wire    [1:0] mm_interconnect_1_sdram_controller_s1_byteenable;               // mm_interconnect_1:SDRAM_Controller_s1_byteenable -> SDRAM_Controller:az_be_n
	wire          mm_interconnect_1_sdram_controller_s1_readdatavalid;            // SDRAM_Controller:za_valid -> mm_interconnect_1:SDRAM_Controller_s1_readdatavalid
	wire          mm_interconnect_1_sdram_controller_s1_write;                    // mm_interconnect_1:SDRAM_Controller_s1_write -> SDRAM_Controller:az_wr_n
	wire   [15:0] mm_interconnect_1_sdram_controller_s1_writedata;                // mm_interconnect_1:SDRAM_Controller_s1_writedata -> SDRAM_Controller:az_data
	wire   [31:0] mm_interconnect_1_avalon_frame_writer_avalon_slave_readdata;    // Avalon_Frame_Writer:S_readdata -> mm_interconnect_1:Avalon_Frame_Writer_avalon_slave_readdata
	wire    [3:0] mm_interconnect_1_avalon_frame_writer_avalon_slave_address;     // mm_interconnect_1:Avalon_Frame_Writer_avalon_slave_address -> Avalon_Frame_Writer:S_address
	wire          mm_interconnect_1_avalon_frame_writer_avalon_slave_read;        // mm_interconnect_1:Avalon_Frame_Writer_avalon_slave_read -> Avalon_Frame_Writer:S_read
	wire          mm_interconnect_1_avalon_frame_writer_avalon_slave_write;       // mm_interconnect_1:Avalon_Frame_Writer_avalon_slave_write -> Avalon_Frame_Writer:S_write
	wire   [31:0] mm_interconnect_1_avalon_frame_writer_avalon_slave_writedata;   // mm_interconnect_1:Avalon_Frame_Writer_avalon_slave_writedata -> Avalon_Frame_Writer:S_writedata
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_awburst;                           // ARM_A9_HPS:h2f_lw_AWBURST -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awburst
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_arlen;                             // ARM_A9_HPS:h2f_lw_ARLEN -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arlen
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_wstrb;                             // ARM_A9_HPS:h2f_lw_WSTRB -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_wstrb
	wire          arm_a9_hps_h2f_lw_axi_master_wready;                            // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_wready -> ARM_A9_HPS:h2f_lw_WREADY
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_rid;                               // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_rid -> ARM_A9_HPS:h2f_lw_RID
	wire          arm_a9_hps_h2f_lw_axi_master_rready;                            // ARM_A9_HPS:h2f_lw_RREADY -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_rready
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_awlen;                             // ARM_A9_HPS:h2f_lw_AWLEN -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awlen
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_wid;                               // ARM_A9_HPS:h2f_lw_WID -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_wid
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_arcache;                           // ARM_A9_HPS:h2f_lw_ARCACHE -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arcache
	wire          arm_a9_hps_h2f_lw_axi_master_wvalid;                            // ARM_A9_HPS:h2f_lw_WVALID -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_wvalid
	wire   [20:0] arm_a9_hps_h2f_lw_axi_master_araddr;                            // ARM_A9_HPS:h2f_lw_ARADDR -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_araddr
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_arprot;                            // ARM_A9_HPS:h2f_lw_ARPROT -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arprot
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_awprot;                            // ARM_A9_HPS:h2f_lw_AWPROT -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awprot
	wire   [31:0] arm_a9_hps_h2f_lw_axi_master_wdata;                             // ARM_A9_HPS:h2f_lw_WDATA -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_wdata
	wire          arm_a9_hps_h2f_lw_axi_master_arvalid;                           // ARM_A9_HPS:h2f_lw_ARVALID -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arvalid
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_awcache;                           // ARM_A9_HPS:h2f_lw_AWCACHE -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awcache
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_arid;                              // ARM_A9_HPS:h2f_lw_ARID -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arid
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_arlock;                            // ARM_A9_HPS:h2f_lw_ARLOCK -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arlock
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_awlock;                            // ARM_A9_HPS:h2f_lw_AWLOCK -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awlock
	wire   [20:0] arm_a9_hps_h2f_lw_axi_master_awaddr;                            // ARM_A9_HPS:h2f_lw_AWADDR -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awaddr
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_bresp;                             // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_bresp -> ARM_A9_HPS:h2f_lw_BRESP
	wire          arm_a9_hps_h2f_lw_axi_master_arready;                           // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arready -> ARM_A9_HPS:h2f_lw_ARREADY
	wire   [31:0] arm_a9_hps_h2f_lw_axi_master_rdata;                             // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_rdata -> ARM_A9_HPS:h2f_lw_RDATA
	wire          arm_a9_hps_h2f_lw_axi_master_awready;                           // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awready -> ARM_A9_HPS:h2f_lw_AWREADY
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_arburst;                           // ARM_A9_HPS:h2f_lw_ARBURST -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arburst
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_arsize;                            // ARM_A9_HPS:h2f_lw_ARSIZE -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_arsize
	wire          arm_a9_hps_h2f_lw_axi_master_bready;                            // ARM_A9_HPS:h2f_lw_BREADY -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_bready
	wire          arm_a9_hps_h2f_lw_axi_master_rlast;                             // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_rlast -> ARM_A9_HPS:h2f_lw_RLAST
	wire          arm_a9_hps_h2f_lw_axi_master_wlast;                             // ARM_A9_HPS:h2f_lw_WLAST -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_wlast
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_rresp;                             // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_rresp -> ARM_A9_HPS:h2f_lw_RRESP
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_awid;                              // ARM_A9_HPS:h2f_lw_AWID -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awid
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_bid;                               // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_bid -> ARM_A9_HPS:h2f_lw_BID
	wire          arm_a9_hps_h2f_lw_axi_master_bvalid;                            // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_bvalid -> ARM_A9_HPS:h2f_lw_BVALID
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_awsize;                            // ARM_A9_HPS:h2f_lw_AWSIZE -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awsize
	wire          arm_a9_hps_h2f_lw_axi_master_awvalid;                           // ARM_A9_HPS:h2f_lw_AWVALID -> mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_awvalid
	wire          arm_a9_hps_h2f_lw_axi_master_rvalid;                            // mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_rvalid -> ARM_A9_HPS:h2f_lw_RVALID
	wire   [31:0] mm_interconnect_2_av_config_avalon_av_config_slave_readdata;    // AV_Config:readdata -> mm_interconnect_2:AV_Config_avalon_av_config_slave_readdata
	wire          mm_interconnect_2_av_config_avalon_av_config_slave_waitrequest; // AV_Config:waitrequest -> mm_interconnect_2:AV_Config_avalon_av_config_slave_waitrequest
	wire    [1:0] mm_interconnect_2_av_config_avalon_av_config_slave_address;     // mm_interconnect_2:AV_Config_avalon_av_config_slave_address -> AV_Config:address
	wire          mm_interconnect_2_av_config_avalon_av_config_slave_read;        // mm_interconnect_2:AV_Config_avalon_av_config_slave_read -> AV_Config:read
	wire    [3:0] mm_interconnect_2_av_config_avalon_av_config_slave_byteenable;  // mm_interconnect_2:AV_Config_avalon_av_config_slave_byteenable -> AV_Config:byteenable
	wire          mm_interconnect_2_av_config_avalon_av_config_slave_write;       // mm_interconnect_2:AV_Config_avalon_av_config_slave_write -> AV_Config:write
	wire   [31:0] mm_interconnect_2_av_config_avalon_av_config_slave_writedata;   // mm_interconnect_2:AV_Config_avalon_av_config_slave_writedata -> AV_Config:writedata
	wire   [31:0] mm_interconnect_2_dot_product_avalon_slave_readdata;            // Dot_Product:slave_readdata -> mm_interconnect_2:Dot_Product_avalon_slave_readdata
	wire          mm_interconnect_2_dot_product_avalon_slave_waitrequest;         // Dot_Product:slave_waitrequest -> mm_interconnect_2:Dot_Product_avalon_slave_waitrequest
	wire    [3:0] mm_interconnect_2_dot_product_avalon_slave_address;             // mm_interconnect_2:Dot_Product_avalon_slave_address -> Dot_Product:slave_address
	wire          mm_interconnect_2_dot_product_avalon_slave_read;                // mm_interconnect_2:Dot_Product_avalon_slave_read -> Dot_Product:slave_read
	wire          mm_interconnect_2_dot_product_avalon_slave_write;               // mm_interconnect_2:Dot_Product_avalon_slave_write -> Dot_Product:slave_write
	wire   [31:0] mm_interconnect_2_dot_product_avalon_slave_writedata;           // mm_interconnect_2:Dot_Product_avalon_slave_writedata -> Dot_Product:slave_writedata
	wire   [31:0] arm_a9_hps_f2h_irq0_irq;                                        // irq_mapper:sender_irq -> ARM_A9_HPS:f2h_irq_p0
	wire   [31:0] arm_a9_hps_f2h_irq1_irq;                                        // irq_mapper_001:sender_irq -> ARM_A9_HPS:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [AV_Config:reset, Avalon_Frame_Writer:reset_n, Dot_Product:rst_n, SDRAM_Controller:reset_n, SRAM1:reset, SRAM2:reset, System_ID:reset_n, mm_interconnect_0:Avalon_Frame_Writer_reset_reset_bridge_in_reset_reset, mm_interconnect_1:Dot_Product_reset_reset_bridge_in_reset_reset, mm_interconnect_2:AV_Config_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire          rst_controller_reset_out_reset_req;                             // rst_controller:reset_req -> [SRAM1:reset_req, SRAM2:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                             // rst_controller_001:reset_out -> [mm_interconnect_0:ARM_A9_HPS_f2h_sdram1_data_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	Computer_System_ARM_A9_HPS #(
		.F2S_Width (3),
		.S2F_Width (3)
	) arm_a9_hps (
		.mem_a                    (memory_mem_a),                                             //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                                            //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                                            //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                                          //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                           //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                                          //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                                         //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                                         //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                                          //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                                       //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                            //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                           //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                                         //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                           //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                                            //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                                         //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),                          //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),                            //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),                            //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),                            //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),                            //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),                            //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),                            //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),                             //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),                          //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),                          //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),                          //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),                            //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),                            //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),                            //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),                              //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),                              //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),                              //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),                              //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),                              //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),                              //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),                              //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),                               //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),                               //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),                              //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),                               //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),                               //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),                               //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),                               //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),                               //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),                               //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),                               //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),                               //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),                               //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),                               //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),                              //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),                              //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),                              //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),                              //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),                             //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),                            //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),                            //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),                             //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),                              //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),                              //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),                              //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),                              //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),                              //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),                              //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),                           //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),                           //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),                           //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_io_hps_io_gpio_inst_GPIO41),                           //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO48  (hps_io_hps_io_gpio_inst_GPIO48),                           //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),                           //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),                           //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),                           //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (h2f_reset_reset_n),                                        //         h2f_reset.reset_n
		.f2h_sdram0_clk           (pixel_clk_clk),                                            //  f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (),                                                         //   f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (),                                                         //                  .burstcount
		.f2h_sdram0_WAITREQUEST   (),                                                         //                  .waitrequest
		.f2h_sdram0_READDATA      (),                                                         //                  .readdata
		.f2h_sdram0_READDATAVALID (),                                                         //                  .readdatavalid
		.f2h_sdram0_READ          (),                                                         //                  .read
		.f2h_sdram0_WRITEDATA     (),                                                         //                  .writedata
		.f2h_sdram0_BYTEENABLE    (),                                                         //                  .byteenable
		.f2h_sdram0_WRITE         (),                                                         //                  .write
		.f2h_sdram1_clk           (pixel_clk_clk),                                            //  f2h_sdram1_clock.clk
		.f2h_sdram1_ADDRESS       (mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_address),     //   f2h_sdram1_data.address
		.f2h_sdram1_BURSTCOUNT    (mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_burstcount),  //                  .burstcount
		.f2h_sdram1_WAITREQUEST   (mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_waitrequest), //                  .waitrequest
		.f2h_sdram1_WRITEDATA     (mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_writedata),   //                  .writedata
		.f2h_sdram1_BYTEENABLE    (mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_byteenable),  //                  .byteenable
		.f2h_sdram1_WRITE         (mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_write),       //                  .write
		.h2f_axi_clk              (pixel_clk_clk),                                            //     h2f_axi_clock.clk
		.h2f_AWID                 (arm_a9_hps_h2f_axi_master_awid),                           //    h2f_axi_master.awid
		.h2f_AWADDR               (arm_a9_hps_h2f_axi_master_awaddr),                         //                  .awaddr
		.h2f_AWLEN                (arm_a9_hps_h2f_axi_master_awlen),                          //                  .awlen
		.h2f_AWSIZE               (arm_a9_hps_h2f_axi_master_awsize),                         //                  .awsize
		.h2f_AWBURST              (arm_a9_hps_h2f_axi_master_awburst),                        //                  .awburst
		.h2f_AWLOCK               (arm_a9_hps_h2f_axi_master_awlock),                         //                  .awlock
		.h2f_AWCACHE              (arm_a9_hps_h2f_axi_master_awcache),                        //                  .awcache
		.h2f_AWPROT               (arm_a9_hps_h2f_axi_master_awprot),                         //                  .awprot
		.h2f_AWVALID              (arm_a9_hps_h2f_axi_master_awvalid),                        //                  .awvalid
		.h2f_AWREADY              (arm_a9_hps_h2f_axi_master_awready),                        //                  .awready
		.h2f_WID                  (arm_a9_hps_h2f_axi_master_wid),                            //                  .wid
		.h2f_WDATA                (arm_a9_hps_h2f_axi_master_wdata),                          //                  .wdata
		.h2f_WSTRB                (arm_a9_hps_h2f_axi_master_wstrb),                          //                  .wstrb
		.h2f_WLAST                (arm_a9_hps_h2f_axi_master_wlast),                          //                  .wlast
		.h2f_WVALID               (arm_a9_hps_h2f_axi_master_wvalid),                         //                  .wvalid
		.h2f_WREADY               (arm_a9_hps_h2f_axi_master_wready),                         //                  .wready
		.h2f_BID                  (arm_a9_hps_h2f_axi_master_bid),                            //                  .bid
		.h2f_BRESP                (arm_a9_hps_h2f_axi_master_bresp),                          //                  .bresp
		.h2f_BVALID               (arm_a9_hps_h2f_axi_master_bvalid),                         //                  .bvalid
		.h2f_BREADY               (arm_a9_hps_h2f_axi_master_bready),                         //                  .bready
		.h2f_ARID                 (arm_a9_hps_h2f_axi_master_arid),                           //                  .arid
		.h2f_ARADDR               (arm_a9_hps_h2f_axi_master_araddr),                         //                  .araddr
		.h2f_ARLEN                (arm_a9_hps_h2f_axi_master_arlen),                          //                  .arlen
		.h2f_ARSIZE               (arm_a9_hps_h2f_axi_master_arsize),                         //                  .arsize
		.h2f_ARBURST              (arm_a9_hps_h2f_axi_master_arburst),                        //                  .arburst
		.h2f_ARLOCK               (arm_a9_hps_h2f_axi_master_arlock),                         //                  .arlock
		.h2f_ARCACHE              (arm_a9_hps_h2f_axi_master_arcache),                        //                  .arcache
		.h2f_ARPROT               (arm_a9_hps_h2f_axi_master_arprot),                         //                  .arprot
		.h2f_ARVALID              (arm_a9_hps_h2f_axi_master_arvalid),                        //                  .arvalid
		.h2f_ARREADY              (arm_a9_hps_h2f_axi_master_arready),                        //                  .arready
		.h2f_RID                  (arm_a9_hps_h2f_axi_master_rid),                            //                  .rid
		.h2f_RDATA                (arm_a9_hps_h2f_axi_master_rdata),                          //                  .rdata
		.h2f_RRESP                (arm_a9_hps_h2f_axi_master_rresp),                          //                  .rresp
		.h2f_RLAST                (arm_a9_hps_h2f_axi_master_rlast),                          //                  .rlast
		.h2f_RVALID               (arm_a9_hps_h2f_axi_master_rvalid),                         //                  .rvalid
		.h2f_RREADY               (arm_a9_hps_h2f_axi_master_rready),                         //                  .rready
		.f2h_axi_clk              (pixel_clk_clk),                                            //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                                         //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                                         //                  .awaddr
		.f2h_AWLEN                (),                                                         //                  .awlen
		.f2h_AWSIZE               (),                                                         //                  .awsize
		.f2h_AWBURST              (),                                                         //                  .awburst
		.f2h_AWLOCK               (),                                                         //                  .awlock
		.f2h_AWCACHE              (),                                                         //                  .awcache
		.f2h_AWPROT               (),                                                         //                  .awprot
		.f2h_AWVALID              (),                                                         //                  .awvalid
		.f2h_AWREADY              (),                                                         //                  .awready
		.f2h_AWUSER               (),                                                         //                  .awuser
		.f2h_WID                  (),                                                         //                  .wid
		.f2h_WDATA                (),                                                         //                  .wdata
		.f2h_WSTRB                (),                                                         //                  .wstrb
		.f2h_WLAST                (),                                                         //                  .wlast
		.f2h_WVALID               (),                                                         //                  .wvalid
		.f2h_WREADY               (),                                                         //                  .wready
		.f2h_BID                  (),                                                         //                  .bid
		.f2h_BRESP                (),                                                         //                  .bresp
		.f2h_BVALID               (),                                                         //                  .bvalid
		.f2h_BREADY               (),                                                         //                  .bready
		.f2h_ARID                 (),                                                         //                  .arid
		.f2h_ARADDR               (),                                                         //                  .araddr
		.f2h_ARLEN                (),                                                         //                  .arlen
		.f2h_ARSIZE               (),                                                         //                  .arsize
		.f2h_ARBURST              (),                                                         //                  .arburst
		.f2h_ARLOCK               (),                                                         //                  .arlock
		.f2h_ARCACHE              (),                                                         //                  .arcache
		.f2h_ARPROT               (),                                                         //                  .arprot
		.f2h_ARVALID              (),                                                         //                  .arvalid
		.f2h_ARREADY              (),                                                         //                  .arready
		.f2h_ARUSER               (),                                                         //                  .aruser
		.f2h_RID                  (),                                                         //                  .rid
		.f2h_RDATA                (),                                                         //                  .rdata
		.f2h_RRESP                (),                                                         //                  .rresp
		.f2h_RLAST                (),                                                         //                  .rlast
		.f2h_RVALID               (),                                                         //                  .rvalid
		.f2h_RREADY               (),                                                         //                  .rready
		.h2f_lw_axi_clk           (pixel_clk_clk),                                            //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (arm_a9_hps_h2f_lw_axi_master_awid),                        // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (arm_a9_hps_h2f_lw_axi_master_awaddr),                      //                  .awaddr
		.h2f_lw_AWLEN             (arm_a9_hps_h2f_lw_axi_master_awlen),                       //                  .awlen
		.h2f_lw_AWSIZE            (arm_a9_hps_h2f_lw_axi_master_awsize),                      //                  .awsize
		.h2f_lw_AWBURST           (arm_a9_hps_h2f_lw_axi_master_awburst),                     //                  .awburst
		.h2f_lw_AWLOCK            (arm_a9_hps_h2f_lw_axi_master_awlock),                      //                  .awlock
		.h2f_lw_AWCACHE           (arm_a9_hps_h2f_lw_axi_master_awcache),                     //                  .awcache
		.h2f_lw_AWPROT            (arm_a9_hps_h2f_lw_axi_master_awprot),                      //                  .awprot
		.h2f_lw_AWVALID           (arm_a9_hps_h2f_lw_axi_master_awvalid),                     //                  .awvalid
		.h2f_lw_AWREADY           (arm_a9_hps_h2f_lw_axi_master_awready),                     //                  .awready
		.h2f_lw_WID               (arm_a9_hps_h2f_lw_axi_master_wid),                         //                  .wid
		.h2f_lw_WDATA             (arm_a9_hps_h2f_lw_axi_master_wdata),                       //                  .wdata
		.h2f_lw_WSTRB             (arm_a9_hps_h2f_lw_axi_master_wstrb),                       //                  .wstrb
		.h2f_lw_WLAST             (arm_a9_hps_h2f_lw_axi_master_wlast),                       //                  .wlast
		.h2f_lw_WVALID            (arm_a9_hps_h2f_lw_axi_master_wvalid),                      //                  .wvalid
		.h2f_lw_WREADY            (arm_a9_hps_h2f_lw_axi_master_wready),                      //                  .wready
		.h2f_lw_BID               (arm_a9_hps_h2f_lw_axi_master_bid),                         //                  .bid
		.h2f_lw_BRESP             (arm_a9_hps_h2f_lw_axi_master_bresp),                       //                  .bresp
		.h2f_lw_BVALID            (arm_a9_hps_h2f_lw_axi_master_bvalid),                      //                  .bvalid
		.h2f_lw_BREADY            (arm_a9_hps_h2f_lw_axi_master_bready),                      //                  .bready
		.h2f_lw_ARID              (arm_a9_hps_h2f_lw_axi_master_arid),                        //                  .arid
		.h2f_lw_ARADDR            (arm_a9_hps_h2f_lw_axi_master_araddr),                      //                  .araddr
		.h2f_lw_ARLEN             (arm_a9_hps_h2f_lw_axi_master_arlen),                       //                  .arlen
		.h2f_lw_ARSIZE            (arm_a9_hps_h2f_lw_axi_master_arsize),                      //                  .arsize
		.h2f_lw_ARBURST           (arm_a9_hps_h2f_lw_axi_master_arburst),                     //                  .arburst
		.h2f_lw_ARLOCK            (arm_a9_hps_h2f_lw_axi_master_arlock),                      //                  .arlock
		.h2f_lw_ARCACHE           (arm_a9_hps_h2f_lw_axi_master_arcache),                     //                  .arcache
		.h2f_lw_ARPROT            (arm_a9_hps_h2f_lw_axi_master_arprot),                      //                  .arprot
		.h2f_lw_ARVALID           (arm_a9_hps_h2f_lw_axi_master_arvalid),                     //                  .arvalid
		.h2f_lw_ARREADY           (arm_a9_hps_h2f_lw_axi_master_arready),                     //                  .arready
		.h2f_lw_RID               (arm_a9_hps_h2f_lw_axi_master_rid),                         //                  .rid
		.h2f_lw_RDATA             (arm_a9_hps_h2f_lw_axi_master_rdata),                       //                  .rdata
		.h2f_lw_RRESP             (arm_a9_hps_h2f_lw_axi_master_rresp),                       //                  .rresp
		.h2f_lw_RLAST             (arm_a9_hps_h2f_lw_axi_master_rlast),                       //                  .rlast
		.h2f_lw_RVALID            (arm_a9_hps_h2f_lw_axi_master_rvalid),                      //                  .rvalid
		.h2f_lw_RREADY            (arm_a9_hps_h2f_lw_axi_master_rready),                      //                  .rready
		.f2h_irq_p0               (arm_a9_hps_f2h_irq0_irq),                                  //          f2h_irq0.irq
		.f2h_irq_p1               (arm_a9_hps_f2h_irq1_irq)                                   //          f2h_irq1.irq
	);

	Computer_System_AV_Config av_config (
		.clk         (pixel_clk_clk),                                                  //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                                 //                  reset.reset
		.address     (mm_interconnect_2_av_config_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_2_av_config_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_2_av_config_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_2_av_config_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_2_av_config_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_2_av_config_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_2_av_config_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (av_config_SDAT),                                                 //     external_interface.export
		.I2C_SCLK    (av_config_SCLK)                                                  //                       .export
	);

	avalon_image_writer #(
		.COMPONENT_SIZE    (8),
		.NUMBER_COMPONENTS (4),
		.PIX_WR            (4)
	) avalon_frame_writer (
		.clk            (pixel_clk_clk),                                                //             clock.clk
		.reset_n        (~rst_controller_reset_out_reset),                              //             reset.reset_n
		.S_address      (mm_interconnect_1_avalon_frame_writer_avalon_slave_address),   //      avalon_slave.address
		.S_writedata    (mm_interconnect_1_avalon_frame_writer_avalon_slave_writedata), //                  .writedata
		.S_readdata     (mm_interconnect_1_avalon_frame_writer_avalon_slave_readdata),  //                  .readdata
		.S_write        (mm_interconnect_1_avalon_frame_writer_avalon_slave_write),     //                  .write
		.S_read         (mm_interconnect_1_avalon_frame_writer_avalon_slave_read),      //                  .read
		.M_address      (avalon_frame_writer_avalon_master_address),                    //     avalon_master.address
		.M_write        (avalon_frame_writer_avalon_master_write),                      //                  .write
		.M_byteenable   (avalon_frame_writer_avalon_master_byteenable),                 //                  .byteenable
		.M_writedata    (avalon_frame_writer_avalon_master_writedata),                  //                  .writedata
		.M_waitrequest  (avalon_frame_writer_avalon_master_waitrequest),                //                  .waitrequest
		.M_burstcount   (avalon_frame_writer_avalon_master_burstcount),                 //                  .burstcount
		.data_valid     (rgba_image_sink_data_valid),                                   //       conduit_end.data_valid
		.input_data     (rgba_image_sink_input_data),                                   //                  .input_data
		.img_width      (rgba_image_sink_img_width),                                    //                  .img_width
		.img_height     (rgba_image_sink_img_height),                                   //                  .img_height
		.stream_reset_n (rgba_stream_reset_reset_n)                                     // stream_reset_sink.reset_n
	);

	dot dot_product (
		.clk                  (pixel_clk_clk),                                          //         clock.clk
		.master_waitrequest   (dot_product_avalon_master_waitrequest),                  // avalon_master.waitrequest
		.master_address       (dot_product_avalon_master_address),                      //              .address
		.master_read          (dot_product_avalon_master_read),                         //              .read
		.master_readdata      (dot_product_avalon_master_readdata),                     //              .readdata
		.master_readdatavalid (dot_product_avalon_master_readdatavalid),                //              .readdatavalid
		.master_write         (dot_product_avalon_master_write),                        //              .write
		.master_writedata     (dot_product_avalon_master_writedata),                    //              .writedata
		.rst_n                (~rst_controller_reset_out_reset),                        //         reset.reset_n
		.slave_waitrequest    (mm_interconnect_2_dot_product_avalon_slave_waitrequest), //  avalon_slave.waitrequest
		.slave_address        (mm_interconnect_2_dot_product_avalon_slave_address),     //              .address
		.slave_read           (mm_interconnect_2_dot_product_avalon_slave_read),        //              .read
		.slave_readdata       (mm_interconnect_2_dot_product_avalon_slave_readdata),    //              .readdata
		.slave_write          (mm_interconnect_2_dot_product_avalon_slave_write),       //              .write
		.slave_writedata      (mm_interconnect_2_dot_product_avalon_slave_writedata)    //              .writedata
	);

	Computer_System_PLL_VGA pll_vga (
		.refclk   (pixel_clk_clk),                 //  refclk.clk
		.rst      (system_pll_reset_source_reset), //   reset.reset
		.outclk_0 (pll_vga_clk_25_clk),            // outclk0.clk
		.locked   ()                               // (terminated)
	);

	Computer_System_SDRAM_Controller sdram_controller (
		.clk            (pixel_clk_clk),                                       //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                     // reset.reset_n
		.az_addr        (mm_interconnect_1_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_1_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_1_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_1_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_1_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_1_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_1_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_1_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_1_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_ctrl_addr),                                     //  wire.export
		.zs_ba          (sdram_ctrl_ba),                                       //      .export
		.zs_cas_n       (sdram_ctrl_cas_n),                                    //      .export
		.zs_cke         (sdram_ctrl_cke),                                      //      .export
		.zs_cs_n        (sdram_ctrl_cs_n),                                     //      .export
		.zs_dq          (sdram_ctrl_dq),                                       //      .export
		.zs_dqm         (sdram_ctrl_dqm),                                      //      .export
		.zs_ras_n       (sdram_ctrl_ras_n),                                    //      .export
		.zs_we_n        (sdram_ctrl_we_n)                                      //      .export
	);

	Computer_System_SRAM1 sram1 (
		.clk        (pixel_clk_clk),                         //   clk1.clk
		.address    (mm_interconnect_1_sram1_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_sram1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_sram1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_sram1_s1_write),      //       .write
		.readdata   (mm_interconnect_1_sram1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_sram1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_sram1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze     (1'b0)                                   // (terminated)
	);

	Computer_System_SRAM2 sram2 (
		.clk        (pixel_clk_clk),                         //   clk1.clk
		.address    (mm_interconnect_1_sram2_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_sram2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_sram2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_sram2_s1_write),      //       .write
		.readdata   (mm_interconnect_1_sram2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_sram2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_sram2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze     (1'b0)                                   // (terminated)
	);

	Computer_System_System_ID system_id (
		.clock    (pixel_clk_clk),                   //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset), //         reset.reset_n
		.readdata (),                                // control_slave.readdata
		.address  ()                                 //              .address
	);

	Computer_System_System_PLL system_pll (
		.ref_clk_clk        (system_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (system_pll_ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (pixel_clk_clk),                 //      sys_clk.clk
		.sdram_clk_clk      (),                              //    sdram_clk.clk
		.reset_source_reset (system_pll_reset_source_reset)  // reset_source.reset
	);

	Computer_System_Video_Subsystem video_subsystem (
		.clk_clk                                                 (pixel_clk_clk),                                                           //                                       clk.clk
		.reset_reset_n                                           (~system_pll_reset_source_reset),                                          //                                     reset.reset_n
		.rgba_image_data                                         (rgba_image_src_data),                                                     //                                rgba_image.data
		.rgba_image_valid                                        (rgba_image_src_valid),                                                    //                                          .valid
		.stream_control_endofpacket                              (stream_control_endofpacket),                                              //                            stream_control.endofpacket
		.stream_control_ready                                    (stream_control_ready),                                                    //                                          .ready
		.stream_control_sreset                                   (stream_control_sreset),                                                   //                                          .sreset
		.video_in_TD_CLK27                                       (video_in_TD_CLK27),                                                       //                                  video_in.TD_CLK27
		.video_in_TD_DATA                                        (video_in_TD_DATA),                                                        //                                          .TD_DATA
		.video_in_TD_HS                                          (video_in_TD_HS),                                                          //                                          .TD_HS
		.video_in_TD_VS                                          (video_in_TD_VS),                                                          //                                          .TD_VS
		.video_in_clk27_reset                                    (video_in_clk27_reset),                                                    //                                          .clk27_reset
		.video_in_TD_RESET                                       (video_in_TD_RESET),                                                       //                                          .TD_RESET
		.video_in_overflow_flag                                  (video_in_overflow_flag),                                                  //                                          .overflow_flag
		.video_in_feed_forward_avalon_forward_sink_data          (video_subsystem_video_in_feed_forward_avalon_forward_sink_data),          // video_in_feed_forward_avalon_forward_sink.data
		.video_in_feed_forward_avalon_forward_sink_startofpacket (video_subsystem_video_in_feed_forward_avalon_forward_sink_startofpacket), //                                          .startofpacket
		.video_in_feed_forward_avalon_forward_sink_endofpacket   (video_subsystem_video_in_feed_forward_avalon_forward_sink_endofpacket),   //                                          .endofpacket
		.video_in_feed_forward_avalon_forward_sink_empty         (video_subsystem_video_in_feed_forward_avalon_forward_sink_empty),         //                                          .empty
		.video_in_feed_forward_avalon_forward_sink_valid         (video_subsystem_video_in_feed_forward_avalon_forward_sink_valid),         //                                          .valid
		.video_in_feed_forward_avalon_forward_sink_ready         (video_subsystem_video_in_feed_forward_avalon_forward_sink_ready),         //                                          .ready
		.video_in_scaler_avalon_scaler_source_ready              (video_subsystem_video_in_scaler_avalon_scaler_source_ready),              //      video_in_scaler_avalon_scaler_source.ready
		.video_in_scaler_avalon_scaler_source_startofpacket      (video_subsystem_video_in_scaler_avalon_scaler_source_startofpacket),      //                                          .startofpacket
		.video_in_scaler_avalon_scaler_source_endofpacket        (video_subsystem_video_in_scaler_avalon_scaler_source_endofpacket),        //                                          .endofpacket
		.video_in_scaler_avalon_scaler_source_valid              (video_subsystem_video_in_scaler_avalon_scaler_source_valid),              //                                          .valid
		.video_in_scaler_avalon_scaler_source_data               (video_subsystem_video_in_scaler_avalon_scaler_source_data)                //                                          .data
	);

	Computer_System_mm_interconnect_0 mm_interconnect_0 (
		.System_PLL_sys_clk_clk                                                  (pixel_clk_clk),                                            //                                                System_PLL_sys_clk.clk
		.ARM_A9_HPS_f2h_sdram1_data_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                       // ARM_A9_HPS_f2h_sdram1_data_translator_reset_reset_bridge_in_reset.reset
		.Avalon_Frame_Writer_reset_reset_bridge_in_reset_reset                   (rst_controller_reset_out_reset),                           //                   Avalon_Frame_Writer_reset_reset_bridge_in_reset.reset
		.Avalon_Frame_Writer_avalon_master_address                               (avalon_frame_writer_avalon_master_address),                //                                 Avalon_Frame_Writer_avalon_master.address
		.Avalon_Frame_Writer_avalon_master_waitrequest                           (avalon_frame_writer_avalon_master_waitrequest),            //                                                                  .waitrequest
		.Avalon_Frame_Writer_avalon_master_burstcount                            (avalon_frame_writer_avalon_master_burstcount),             //                                                                  .burstcount
		.Avalon_Frame_Writer_avalon_master_byteenable                            (avalon_frame_writer_avalon_master_byteenable),             //                                                                  .byteenable
		.Avalon_Frame_Writer_avalon_master_write                                 (avalon_frame_writer_avalon_master_write),                  //                                                                  .write
		.Avalon_Frame_Writer_avalon_master_writedata                             (avalon_frame_writer_avalon_master_writedata),              //                                                                  .writedata
		.ARM_A9_HPS_f2h_sdram1_data_address                                      (mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_address),     //                                        ARM_A9_HPS_f2h_sdram1_data.address
		.ARM_A9_HPS_f2h_sdram1_data_write                                        (mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_write),       //                                                                  .write
		.ARM_A9_HPS_f2h_sdram1_data_writedata                                    (mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_writedata),   //                                                                  .writedata
		.ARM_A9_HPS_f2h_sdram1_data_burstcount                                   (mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_burstcount),  //                                                                  .burstcount
		.ARM_A9_HPS_f2h_sdram1_data_byteenable                                   (mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_byteenable),  //                                                                  .byteenable
		.ARM_A9_HPS_f2h_sdram1_data_waitrequest                                  (mm_interconnect_0_arm_a9_hps_f2h_sdram1_data_waitrequest)  //                                                                  .waitrequest
	);

	Computer_System_mm_interconnect_1 mm_interconnect_1 (
		.ARM_A9_HPS_h2f_axi_master_awid                                        (arm_a9_hps_h2f_axi_master_awid),                               //                                       ARM_A9_HPS_h2f_axi_master.awid
		.ARM_A9_HPS_h2f_axi_master_awaddr                                      (arm_a9_hps_h2f_axi_master_awaddr),                             //                                                                .awaddr
		.ARM_A9_HPS_h2f_axi_master_awlen                                       (arm_a9_hps_h2f_axi_master_awlen),                              //                                                                .awlen
		.ARM_A9_HPS_h2f_axi_master_awsize                                      (arm_a9_hps_h2f_axi_master_awsize),                             //                                                                .awsize
		.ARM_A9_HPS_h2f_axi_master_awburst                                     (arm_a9_hps_h2f_axi_master_awburst),                            //                                                                .awburst
		.ARM_A9_HPS_h2f_axi_master_awlock                                      (arm_a9_hps_h2f_axi_master_awlock),                             //                                                                .awlock
		.ARM_A9_HPS_h2f_axi_master_awcache                                     (arm_a9_hps_h2f_axi_master_awcache),                            //                                                                .awcache
		.ARM_A9_HPS_h2f_axi_master_awprot                                      (arm_a9_hps_h2f_axi_master_awprot),                             //                                                                .awprot
		.ARM_A9_HPS_h2f_axi_master_awvalid                                     (arm_a9_hps_h2f_axi_master_awvalid),                            //                                                                .awvalid
		.ARM_A9_HPS_h2f_axi_master_awready                                     (arm_a9_hps_h2f_axi_master_awready),                            //                                                                .awready
		.ARM_A9_HPS_h2f_axi_master_wid                                         (arm_a9_hps_h2f_axi_master_wid),                                //                                                                .wid
		.ARM_A9_HPS_h2f_axi_master_wdata                                       (arm_a9_hps_h2f_axi_master_wdata),                              //                                                                .wdata
		.ARM_A9_HPS_h2f_axi_master_wstrb                                       (arm_a9_hps_h2f_axi_master_wstrb),                              //                                                                .wstrb
		.ARM_A9_HPS_h2f_axi_master_wlast                                       (arm_a9_hps_h2f_axi_master_wlast),                              //                                                                .wlast
		.ARM_A9_HPS_h2f_axi_master_wvalid                                      (arm_a9_hps_h2f_axi_master_wvalid),                             //                                                                .wvalid
		.ARM_A9_HPS_h2f_axi_master_wready                                      (arm_a9_hps_h2f_axi_master_wready),                             //                                                                .wready
		.ARM_A9_HPS_h2f_axi_master_bid                                         (arm_a9_hps_h2f_axi_master_bid),                                //                                                                .bid
		.ARM_A9_HPS_h2f_axi_master_bresp                                       (arm_a9_hps_h2f_axi_master_bresp),                              //                                                                .bresp
		.ARM_A9_HPS_h2f_axi_master_bvalid                                      (arm_a9_hps_h2f_axi_master_bvalid),                             //                                                                .bvalid
		.ARM_A9_HPS_h2f_axi_master_bready                                      (arm_a9_hps_h2f_axi_master_bready),                             //                                                                .bready
		.ARM_A9_HPS_h2f_axi_master_arid                                        (arm_a9_hps_h2f_axi_master_arid),                               //                                                                .arid
		.ARM_A9_HPS_h2f_axi_master_araddr                                      (arm_a9_hps_h2f_axi_master_araddr),                             //                                                                .araddr
		.ARM_A9_HPS_h2f_axi_master_arlen                                       (arm_a9_hps_h2f_axi_master_arlen),                              //                                                                .arlen
		.ARM_A9_HPS_h2f_axi_master_arsize                                      (arm_a9_hps_h2f_axi_master_arsize),                             //                                                                .arsize
		.ARM_A9_HPS_h2f_axi_master_arburst                                     (arm_a9_hps_h2f_axi_master_arburst),                            //                                                                .arburst
		.ARM_A9_HPS_h2f_axi_master_arlock                                      (arm_a9_hps_h2f_axi_master_arlock),                             //                                                                .arlock
		.ARM_A9_HPS_h2f_axi_master_arcache                                     (arm_a9_hps_h2f_axi_master_arcache),                            //                                                                .arcache
		.ARM_A9_HPS_h2f_axi_master_arprot                                      (arm_a9_hps_h2f_axi_master_arprot),                             //                                                                .arprot
		.ARM_A9_HPS_h2f_axi_master_arvalid                                     (arm_a9_hps_h2f_axi_master_arvalid),                            //                                                                .arvalid
		.ARM_A9_HPS_h2f_axi_master_arready                                     (arm_a9_hps_h2f_axi_master_arready),                            //                                                                .arready
		.ARM_A9_HPS_h2f_axi_master_rid                                         (arm_a9_hps_h2f_axi_master_rid),                                //                                                                .rid
		.ARM_A9_HPS_h2f_axi_master_rdata                                       (arm_a9_hps_h2f_axi_master_rdata),                              //                                                                .rdata
		.ARM_A9_HPS_h2f_axi_master_rresp                                       (arm_a9_hps_h2f_axi_master_rresp),                              //                                                                .rresp
		.ARM_A9_HPS_h2f_axi_master_rlast                                       (arm_a9_hps_h2f_axi_master_rlast),                              //                                                                .rlast
		.ARM_A9_HPS_h2f_axi_master_rvalid                                      (arm_a9_hps_h2f_axi_master_rvalid),                             //                                                                .rvalid
		.ARM_A9_HPS_h2f_axi_master_rready                                      (arm_a9_hps_h2f_axi_master_rready),                             //                                                                .rready
		.System_PLL_sys_clk_clk                                                (pixel_clk_clk),                                                //                                              System_PLL_sys_clk.clk
		.ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                           // ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.Dot_Product_reset_reset_bridge_in_reset_reset                         (rst_controller_reset_out_reset),                               //                         Dot_Product_reset_reset_bridge_in_reset.reset
		.Dot_Product_avalon_master_address                                     (dot_product_avalon_master_address),                            //                                       Dot_Product_avalon_master.address
		.Dot_Product_avalon_master_waitrequest                                 (dot_product_avalon_master_waitrequest),                        //                                                                .waitrequest
		.Dot_Product_avalon_master_read                                        (dot_product_avalon_master_read),                               //                                                                .read
		.Dot_Product_avalon_master_readdata                                    (dot_product_avalon_master_readdata),                           //                                                                .readdata
		.Dot_Product_avalon_master_readdatavalid                               (dot_product_avalon_master_readdatavalid),                      //                                                                .readdatavalid
		.Dot_Product_avalon_master_write                                       (dot_product_avalon_master_write),                              //                                                                .write
		.Dot_Product_avalon_master_writedata                                   (dot_product_avalon_master_writedata),                          //                                                                .writedata
		.Avalon_Frame_Writer_avalon_slave_address                              (mm_interconnect_1_avalon_frame_writer_avalon_slave_address),   //                                Avalon_Frame_Writer_avalon_slave.address
		.Avalon_Frame_Writer_avalon_slave_write                                (mm_interconnect_1_avalon_frame_writer_avalon_slave_write),     //                                                                .write
		.Avalon_Frame_Writer_avalon_slave_read                                 (mm_interconnect_1_avalon_frame_writer_avalon_slave_read),      //                                                                .read
		.Avalon_Frame_Writer_avalon_slave_readdata                             (mm_interconnect_1_avalon_frame_writer_avalon_slave_readdata),  //                                                                .readdata
		.Avalon_Frame_Writer_avalon_slave_writedata                            (mm_interconnect_1_avalon_frame_writer_avalon_slave_writedata), //                                                                .writedata
		.SDRAM_Controller_s1_address                                           (mm_interconnect_1_sdram_controller_s1_address),                //                                             SDRAM_Controller_s1.address
		.SDRAM_Controller_s1_write                                             (mm_interconnect_1_sdram_controller_s1_write),                  //                                                                .write
		.SDRAM_Controller_s1_read                                              (mm_interconnect_1_sdram_controller_s1_read),                   //                                                                .read
		.SDRAM_Controller_s1_readdata                                          (mm_interconnect_1_sdram_controller_s1_readdata),               //                                                                .readdata
		.SDRAM_Controller_s1_writedata                                         (mm_interconnect_1_sdram_controller_s1_writedata),              //                                                                .writedata
		.SDRAM_Controller_s1_byteenable                                        (mm_interconnect_1_sdram_controller_s1_byteenable),             //                                                                .byteenable
		.SDRAM_Controller_s1_readdatavalid                                     (mm_interconnect_1_sdram_controller_s1_readdatavalid),          //                                                                .readdatavalid
		.SDRAM_Controller_s1_waitrequest                                       (mm_interconnect_1_sdram_controller_s1_waitrequest),            //                                                                .waitrequest
		.SDRAM_Controller_s1_chipselect                                        (mm_interconnect_1_sdram_controller_s1_chipselect),             //                                                                .chipselect
		.SRAM1_s1_address                                                      (mm_interconnect_1_sram1_s1_address),                           //                                                        SRAM1_s1.address
		.SRAM1_s1_write                                                        (mm_interconnect_1_sram1_s1_write),                             //                                                                .write
		.SRAM1_s1_readdata                                                     (mm_interconnect_1_sram1_s1_readdata),                          //                                                                .readdata
		.SRAM1_s1_writedata                                                    (mm_interconnect_1_sram1_s1_writedata),                         //                                                                .writedata
		.SRAM1_s1_byteenable                                                   (mm_interconnect_1_sram1_s1_byteenable),                        //                                                                .byteenable
		.SRAM1_s1_chipselect                                                   (mm_interconnect_1_sram1_s1_chipselect),                        //                                                                .chipselect
		.SRAM1_s1_clken                                                        (mm_interconnect_1_sram1_s1_clken),                             //                                                                .clken
		.SRAM2_s1_address                                                      (mm_interconnect_1_sram2_s1_address),                           //                                                        SRAM2_s1.address
		.SRAM2_s1_write                                                        (mm_interconnect_1_sram2_s1_write),                             //                                                                .write
		.SRAM2_s1_readdata                                                     (mm_interconnect_1_sram2_s1_readdata),                          //                                                                .readdata
		.SRAM2_s1_writedata                                                    (mm_interconnect_1_sram2_s1_writedata),                         //                                                                .writedata
		.SRAM2_s1_byteenable                                                   (mm_interconnect_1_sram2_s1_byteenable),                        //                                                                .byteenable
		.SRAM2_s1_chipselect                                                   (mm_interconnect_1_sram2_s1_chipselect),                        //                                                                .chipselect
		.SRAM2_s1_clken                                                        (mm_interconnect_1_sram2_s1_clken)                              //                                                                .clken
	);

	Computer_System_mm_interconnect_2 mm_interconnect_2 (
		.ARM_A9_HPS_h2f_lw_axi_master_awid                                        (arm_a9_hps_h2f_lw_axi_master_awid),                              //                                       ARM_A9_HPS_h2f_lw_axi_master.awid
		.ARM_A9_HPS_h2f_lw_axi_master_awaddr                                      (arm_a9_hps_h2f_lw_axi_master_awaddr),                            //                                                                   .awaddr
		.ARM_A9_HPS_h2f_lw_axi_master_awlen                                       (arm_a9_hps_h2f_lw_axi_master_awlen),                             //                                                                   .awlen
		.ARM_A9_HPS_h2f_lw_axi_master_awsize                                      (arm_a9_hps_h2f_lw_axi_master_awsize),                            //                                                                   .awsize
		.ARM_A9_HPS_h2f_lw_axi_master_awburst                                     (arm_a9_hps_h2f_lw_axi_master_awburst),                           //                                                                   .awburst
		.ARM_A9_HPS_h2f_lw_axi_master_awlock                                      (arm_a9_hps_h2f_lw_axi_master_awlock),                            //                                                                   .awlock
		.ARM_A9_HPS_h2f_lw_axi_master_awcache                                     (arm_a9_hps_h2f_lw_axi_master_awcache),                           //                                                                   .awcache
		.ARM_A9_HPS_h2f_lw_axi_master_awprot                                      (arm_a9_hps_h2f_lw_axi_master_awprot),                            //                                                                   .awprot
		.ARM_A9_HPS_h2f_lw_axi_master_awvalid                                     (arm_a9_hps_h2f_lw_axi_master_awvalid),                           //                                                                   .awvalid
		.ARM_A9_HPS_h2f_lw_axi_master_awready                                     (arm_a9_hps_h2f_lw_axi_master_awready),                           //                                                                   .awready
		.ARM_A9_HPS_h2f_lw_axi_master_wid                                         (arm_a9_hps_h2f_lw_axi_master_wid),                               //                                                                   .wid
		.ARM_A9_HPS_h2f_lw_axi_master_wdata                                       (arm_a9_hps_h2f_lw_axi_master_wdata),                             //                                                                   .wdata
		.ARM_A9_HPS_h2f_lw_axi_master_wstrb                                       (arm_a9_hps_h2f_lw_axi_master_wstrb),                             //                                                                   .wstrb
		.ARM_A9_HPS_h2f_lw_axi_master_wlast                                       (arm_a9_hps_h2f_lw_axi_master_wlast),                             //                                                                   .wlast
		.ARM_A9_HPS_h2f_lw_axi_master_wvalid                                      (arm_a9_hps_h2f_lw_axi_master_wvalid),                            //                                                                   .wvalid
		.ARM_A9_HPS_h2f_lw_axi_master_wready                                      (arm_a9_hps_h2f_lw_axi_master_wready),                            //                                                                   .wready
		.ARM_A9_HPS_h2f_lw_axi_master_bid                                         (arm_a9_hps_h2f_lw_axi_master_bid),                               //                                                                   .bid
		.ARM_A9_HPS_h2f_lw_axi_master_bresp                                       (arm_a9_hps_h2f_lw_axi_master_bresp),                             //                                                                   .bresp
		.ARM_A9_HPS_h2f_lw_axi_master_bvalid                                      (arm_a9_hps_h2f_lw_axi_master_bvalid),                            //                                                                   .bvalid
		.ARM_A9_HPS_h2f_lw_axi_master_bready                                      (arm_a9_hps_h2f_lw_axi_master_bready),                            //                                                                   .bready
		.ARM_A9_HPS_h2f_lw_axi_master_arid                                        (arm_a9_hps_h2f_lw_axi_master_arid),                              //                                                                   .arid
		.ARM_A9_HPS_h2f_lw_axi_master_araddr                                      (arm_a9_hps_h2f_lw_axi_master_araddr),                            //                                                                   .araddr
		.ARM_A9_HPS_h2f_lw_axi_master_arlen                                       (arm_a9_hps_h2f_lw_axi_master_arlen),                             //                                                                   .arlen
		.ARM_A9_HPS_h2f_lw_axi_master_arsize                                      (arm_a9_hps_h2f_lw_axi_master_arsize),                            //                                                                   .arsize
		.ARM_A9_HPS_h2f_lw_axi_master_arburst                                     (arm_a9_hps_h2f_lw_axi_master_arburst),                           //                                                                   .arburst
		.ARM_A9_HPS_h2f_lw_axi_master_arlock                                      (arm_a9_hps_h2f_lw_axi_master_arlock),                            //                                                                   .arlock
		.ARM_A9_HPS_h2f_lw_axi_master_arcache                                     (arm_a9_hps_h2f_lw_axi_master_arcache),                           //                                                                   .arcache
		.ARM_A9_HPS_h2f_lw_axi_master_arprot                                      (arm_a9_hps_h2f_lw_axi_master_arprot),                            //                                                                   .arprot
		.ARM_A9_HPS_h2f_lw_axi_master_arvalid                                     (arm_a9_hps_h2f_lw_axi_master_arvalid),                           //                                                                   .arvalid
		.ARM_A9_HPS_h2f_lw_axi_master_arready                                     (arm_a9_hps_h2f_lw_axi_master_arready),                           //                                                                   .arready
		.ARM_A9_HPS_h2f_lw_axi_master_rid                                         (arm_a9_hps_h2f_lw_axi_master_rid),                               //                                                                   .rid
		.ARM_A9_HPS_h2f_lw_axi_master_rdata                                       (arm_a9_hps_h2f_lw_axi_master_rdata),                             //                                                                   .rdata
		.ARM_A9_HPS_h2f_lw_axi_master_rresp                                       (arm_a9_hps_h2f_lw_axi_master_rresp),                             //                                                                   .rresp
		.ARM_A9_HPS_h2f_lw_axi_master_rlast                                       (arm_a9_hps_h2f_lw_axi_master_rlast),                             //                                                                   .rlast
		.ARM_A9_HPS_h2f_lw_axi_master_rvalid                                      (arm_a9_hps_h2f_lw_axi_master_rvalid),                            //                                                                   .rvalid
		.ARM_A9_HPS_h2f_lw_axi_master_rready                                      (arm_a9_hps_h2f_lw_axi_master_rready),                            //                                                                   .rready
		.System_PLL_sys_clk_clk                                                   (pixel_clk_clk),                                                  //                                                 System_PLL_sys_clk.clk
		.ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                             // ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.AV_Config_reset_reset_bridge_in_reset_reset                              (rst_controller_reset_out_reset),                                 //                              AV_Config_reset_reset_bridge_in_reset.reset
		.AV_Config_avalon_av_config_slave_address                                 (mm_interconnect_2_av_config_avalon_av_config_slave_address),     //                                   AV_Config_avalon_av_config_slave.address
		.AV_Config_avalon_av_config_slave_write                                   (mm_interconnect_2_av_config_avalon_av_config_slave_write),       //                                                                   .write
		.AV_Config_avalon_av_config_slave_read                                    (mm_interconnect_2_av_config_avalon_av_config_slave_read),        //                                                                   .read
		.AV_Config_avalon_av_config_slave_readdata                                (mm_interconnect_2_av_config_avalon_av_config_slave_readdata),    //                                                                   .readdata
		.AV_Config_avalon_av_config_slave_writedata                               (mm_interconnect_2_av_config_avalon_av_config_slave_writedata),   //                                                                   .writedata
		.AV_Config_avalon_av_config_slave_byteenable                              (mm_interconnect_2_av_config_avalon_av_config_slave_byteenable),  //                                                                   .byteenable
		.AV_Config_avalon_av_config_slave_waitrequest                             (mm_interconnect_2_av_config_avalon_av_config_slave_waitrequest), //                                                                   .waitrequest
		.Dot_Product_avalon_slave_address                                         (mm_interconnect_2_dot_product_avalon_slave_address),             //                                           Dot_Product_avalon_slave.address
		.Dot_Product_avalon_slave_write                                           (mm_interconnect_2_dot_product_avalon_slave_write),               //                                                                   .write
		.Dot_Product_avalon_slave_read                                            (mm_interconnect_2_dot_product_avalon_slave_read),                //                                                                   .read
		.Dot_Product_avalon_slave_readdata                                        (mm_interconnect_2_dot_product_avalon_slave_readdata),            //                                                                   .readdata
		.Dot_Product_avalon_slave_writedata                                       (mm_interconnect_2_dot_product_avalon_slave_writedata),           //                                                                   .writedata
		.Dot_Product_avalon_slave_waitrequest                                     (mm_interconnect_2_dot_product_avalon_slave_waitrequest)          //                                                                   .waitrequest
	);

	Computer_System_irq_mapper irq_mapper (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq0_irq)  //    sender.irq
	);

	Computer_System_irq_mapper irq_mapper_001 (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (system_pll_reset_source_reset),      // reset_in0.reset
		.clk            (pixel_clk_clk),                      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~h2f_reset_reset_n),                 // reset_in0.reset
		.clk            (pixel_clk_clk),                      //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
