
module Computer_System (
	av_config_SDAT,
	av_config_SCLK,
	h2f_reset_reset_n,
	hps_io_hps_io_emac1_inst_TX_CLK,
	hps_io_hps_io_emac1_inst_TXD0,
	hps_io_hps_io_emac1_inst_TXD1,
	hps_io_hps_io_emac1_inst_TXD2,
	hps_io_hps_io_emac1_inst_TXD3,
	hps_io_hps_io_emac1_inst_RXD0,
	hps_io_hps_io_emac1_inst_MDIO,
	hps_io_hps_io_emac1_inst_MDC,
	hps_io_hps_io_emac1_inst_RX_CTL,
	hps_io_hps_io_emac1_inst_TX_CTL,
	hps_io_hps_io_emac1_inst_RX_CLK,
	hps_io_hps_io_emac1_inst_RXD1,
	hps_io_hps_io_emac1_inst_RXD2,
	hps_io_hps_io_emac1_inst_RXD3,
	hps_io_hps_io_qspi_inst_IO0,
	hps_io_hps_io_qspi_inst_IO1,
	hps_io_hps_io_qspi_inst_IO2,
	hps_io_hps_io_qspi_inst_IO3,
	hps_io_hps_io_qspi_inst_SS0,
	hps_io_hps_io_qspi_inst_CLK,
	hps_io_hps_io_sdio_inst_CMD,
	hps_io_hps_io_sdio_inst_D0,
	hps_io_hps_io_sdio_inst_D1,
	hps_io_hps_io_sdio_inst_CLK,
	hps_io_hps_io_sdio_inst_D2,
	hps_io_hps_io_sdio_inst_D3,
	hps_io_hps_io_usb1_inst_D0,
	hps_io_hps_io_usb1_inst_D1,
	hps_io_hps_io_usb1_inst_D2,
	hps_io_hps_io_usb1_inst_D3,
	hps_io_hps_io_usb1_inst_D4,
	hps_io_hps_io_usb1_inst_D5,
	hps_io_hps_io_usb1_inst_D6,
	hps_io_hps_io_usb1_inst_D7,
	hps_io_hps_io_usb1_inst_CLK,
	hps_io_hps_io_usb1_inst_STP,
	hps_io_hps_io_usb1_inst_DIR,
	hps_io_hps_io_usb1_inst_NXT,
	hps_io_hps_io_spim1_inst_CLK,
	hps_io_hps_io_spim1_inst_MOSI,
	hps_io_hps_io_spim1_inst_MISO,
	hps_io_hps_io_spim1_inst_SS0,
	hps_io_hps_io_uart0_inst_RX,
	hps_io_hps_io_uart0_inst_TX,
	hps_io_hps_io_i2c0_inst_SDA,
	hps_io_hps_io_i2c0_inst_SCL,
	hps_io_hps_io_i2c1_inst_SDA,
	hps_io_hps_io_i2c1_inst_SCL,
	hps_io_hps_io_gpio_inst_GPIO09,
	hps_io_hps_io_gpio_inst_GPIO35,
	hps_io_hps_io_gpio_inst_GPIO40,
	hps_io_hps_io_gpio_inst_GPIO41,
	hps_io_hps_io_gpio_inst_GPIO48,
	hps_io_hps_io_gpio_inst_GPIO53,
	hps_io_hps_io_gpio_inst_GPIO54,
	hps_io_hps_io_gpio_inst_GPIO61,
	memory_mem_a,
	memory_mem_ba,
	memory_mem_ck,
	memory_mem_ck_n,
	memory_mem_cke,
	memory_mem_cs_n,
	memory_mem_ras_n,
	memory_mem_cas_n,
	memory_mem_we_n,
	memory_mem_reset_n,
	memory_mem_dq,
	memory_mem_dqs,
	memory_mem_dqs_n,
	memory_mem_odt,
	memory_mem_dm,
	memory_oct_rzqin,
	pixel_clk_clk,
	pll_vga_clk_25_clk,
	rgba_image_sink_data_valid,
	rgba_image_sink_input_data,
	rgba_image_sink_img_width,
	rgba_image_sink_img_height,
	rgba_image_src_data,
	rgba_image_src_valid,
	rgba_stream_reset_reset_n,
	sdram_ctrl_addr,
	sdram_ctrl_ba,
	sdram_ctrl_cas_n,
	sdram_ctrl_cke,
	sdram_ctrl_cs_n,
	sdram_ctrl_dq,
	sdram_ctrl_dqm,
	sdram_ctrl_ras_n,
	sdram_ctrl_we_n,
	stream_control_endofpacket,
	stream_control_ready,
	stream_control_sreset,
	stream_control_startofpacket,
	stream_control_frame_transition,
	system_pll_ref_clk_clk,
	system_pll_ref_reset_reset,
	video_in_TD_CLK27,
	video_in_TD_DATA,
	video_in_TD_HS,
	video_in_TD_VS,
	video_in_clk27_reset,
	video_in_TD_RESET,
	video_in_overflow_flag,
	video_subsystem_video_in_feed_forward_avalon_forward_sink_data,
	video_subsystem_video_in_feed_forward_avalon_forward_sink_startofpacket,
	video_subsystem_video_in_feed_forward_avalon_forward_sink_endofpacket,
	video_subsystem_video_in_feed_forward_avalon_forward_sink_empty,
	video_subsystem_video_in_feed_forward_avalon_forward_sink_valid,
	video_subsystem_video_in_feed_forward_avalon_forward_sink_ready,
	video_subsystem_video_in_scaler_avalon_scaler_source_ready,
	video_subsystem_video_in_scaler_avalon_scaler_source_startofpacket,
	video_subsystem_video_in_scaler_avalon_scaler_source_endofpacket,
	video_subsystem_video_in_scaler_avalon_scaler_source_valid,
	video_subsystem_video_in_scaler_avalon_scaler_source_data,
	video_subsystem_video_in_scaler_avalon_scaler_source_channel);	

	inout		av_config_SDAT;
	output		av_config_SCLK;
	output		h2f_reset_reset_n;
	output		hps_io_hps_io_emac1_inst_TX_CLK;
	output		hps_io_hps_io_emac1_inst_TXD0;
	output		hps_io_hps_io_emac1_inst_TXD1;
	output		hps_io_hps_io_emac1_inst_TXD2;
	output		hps_io_hps_io_emac1_inst_TXD3;
	input		hps_io_hps_io_emac1_inst_RXD0;
	inout		hps_io_hps_io_emac1_inst_MDIO;
	output		hps_io_hps_io_emac1_inst_MDC;
	input		hps_io_hps_io_emac1_inst_RX_CTL;
	output		hps_io_hps_io_emac1_inst_TX_CTL;
	input		hps_io_hps_io_emac1_inst_RX_CLK;
	input		hps_io_hps_io_emac1_inst_RXD1;
	input		hps_io_hps_io_emac1_inst_RXD2;
	input		hps_io_hps_io_emac1_inst_RXD3;
	inout		hps_io_hps_io_qspi_inst_IO0;
	inout		hps_io_hps_io_qspi_inst_IO1;
	inout		hps_io_hps_io_qspi_inst_IO2;
	inout		hps_io_hps_io_qspi_inst_IO3;
	output		hps_io_hps_io_qspi_inst_SS0;
	output		hps_io_hps_io_qspi_inst_CLK;
	inout		hps_io_hps_io_sdio_inst_CMD;
	inout		hps_io_hps_io_sdio_inst_D0;
	inout		hps_io_hps_io_sdio_inst_D1;
	output		hps_io_hps_io_sdio_inst_CLK;
	inout		hps_io_hps_io_sdio_inst_D2;
	inout		hps_io_hps_io_sdio_inst_D3;
	inout		hps_io_hps_io_usb1_inst_D0;
	inout		hps_io_hps_io_usb1_inst_D1;
	inout		hps_io_hps_io_usb1_inst_D2;
	inout		hps_io_hps_io_usb1_inst_D3;
	inout		hps_io_hps_io_usb1_inst_D4;
	inout		hps_io_hps_io_usb1_inst_D5;
	inout		hps_io_hps_io_usb1_inst_D6;
	inout		hps_io_hps_io_usb1_inst_D7;
	input		hps_io_hps_io_usb1_inst_CLK;
	output		hps_io_hps_io_usb1_inst_STP;
	input		hps_io_hps_io_usb1_inst_DIR;
	input		hps_io_hps_io_usb1_inst_NXT;
	output		hps_io_hps_io_spim1_inst_CLK;
	output		hps_io_hps_io_spim1_inst_MOSI;
	input		hps_io_hps_io_spim1_inst_MISO;
	output		hps_io_hps_io_spim1_inst_SS0;
	input		hps_io_hps_io_uart0_inst_RX;
	output		hps_io_hps_io_uart0_inst_TX;
	inout		hps_io_hps_io_i2c0_inst_SDA;
	inout		hps_io_hps_io_i2c0_inst_SCL;
	inout		hps_io_hps_io_i2c1_inst_SDA;
	inout		hps_io_hps_io_i2c1_inst_SCL;
	inout		hps_io_hps_io_gpio_inst_GPIO09;
	inout		hps_io_hps_io_gpio_inst_GPIO35;
	inout		hps_io_hps_io_gpio_inst_GPIO40;
	inout		hps_io_hps_io_gpio_inst_GPIO41;
	inout		hps_io_hps_io_gpio_inst_GPIO48;
	inout		hps_io_hps_io_gpio_inst_GPIO53;
	inout		hps_io_hps_io_gpio_inst_GPIO54;
	inout		hps_io_hps_io_gpio_inst_GPIO61;
	output	[14:0]	memory_mem_a;
	output	[2:0]	memory_mem_ba;
	output		memory_mem_ck;
	output		memory_mem_ck_n;
	output		memory_mem_cke;
	output		memory_mem_cs_n;
	output		memory_mem_ras_n;
	output		memory_mem_cas_n;
	output		memory_mem_we_n;
	output		memory_mem_reset_n;
	inout	[31:0]	memory_mem_dq;
	inout	[3:0]	memory_mem_dqs;
	inout	[3:0]	memory_mem_dqs_n;
	output		memory_mem_odt;
	output	[3:0]	memory_mem_dm;
	input		memory_oct_rzqin;
	output		pixel_clk_clk;
	output		pll_vga_clk_25_clk;
	input		rgba_image_sink_data_valid;
	input	[31:0]	rgba_image_sink_input_data;
	input	[15:0]	rgba_image_sink_img_width;
	input	[15:0]	rgba_image_sink_img_height;
	output	[31:0]	rgba_image_src_data;
	output		rgba_image_src_valid;
	input		rgba_stream_reset_reset_n;
	output	[12:0]	sdram_ctrl_addr;
	output	[1:0]	sdram_ctrl_ba;
	output		sdram_ctrl_cas_n;
	output		sdram_ctrl_cke;
	output		sdram_ctrl_cs_n;
	inout	[15:0]	sdram_ctrl_dq;
	output	[1:0]	sdram_ctrl_dqm;
	output		sdram_ctrl_ras_n;
	output		sdram_ctrl_we_n;
	input		stream_control_endofpacket;
	output		stream_control_ready;
	output		stream_control_sreset;
	input		stream_control_startofpacket;
	output		stream_control_frame_transition;
	input		system_pll_ref_clk_clk;
	input		system_pll_ref_reset_reset;
	input		video_in_TD_CLK27;
	input	[7:0]	video_in_TD_DATA;
	input		video_in_TD_HS;
	input		video_in_TD_VS;
	input		video_in_clk27_reset;
	output		video_in_TD_RESET;
	output		video_in_overflow_flag;
	input	[23:0]	video_subsystem_video_in_feed_forward_avalon_forward_sink_data;
	input		video_subsystem_video_in_feed_forward_avalon_forward_sink_startofpacket;
	input		video_subsystem_video_in_feed_forward_avalon_forward_sink_endofpacket;
	input	[1:0]	video_subsystem_video_in_feed_forward_avalon_forward_sink_empty;
	input		video_subsystem_video_in_feed_forward_avalon_forward_sink_valid;
	output		video_subsystem_video_in_feed_forward_avalon_forward_sink_ready;
	input		video_subsystem_video_in_scaler_avalon_scaler_source_ready;
	output		video_subsystem_video_in_scaler_avalon_scaler_source_startofpacket;
	output		video_subsystem_video_in_scaler_avalon_scaler_source_endofpacket;
	output		video_subsystem_video_in_scaler_avalon_scaler_source_valid;
	output	[23:0]	video_subsystem_video_in_scaler_avalon_scaler_source_data;
	output		video_subsystem_video_in_scaler_avalon_scaler_source_channel;
endmodule
