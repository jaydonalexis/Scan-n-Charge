	component Computer_System is
		port (
			av_config_SDAT                                                          : inout std_logic                     := 'X';             -- SDAT
			av_config_SCLK                                                          : out   std_logic;                                        -- SCLK
			h2f_reset_reset_n                                                       : out   std_logic;                                        -- reset_n
			hps_io_hps_io_emac1_inst_TX_CLK                                         : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_io_hps_io_emac1_inst_TXD0                                           : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_io_hps_io_emac1_inst_TXD1                                           : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_io_hps_io_emac1_inst_TXD2                                           : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_io_hps_io_emac1_inst_TXD3                                           : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_io_hps_io_emac1_inst_RXD0                                           : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_hps_io_emac1_inst_MDIO                                           : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_hps_io_emac1_inst_MDC                                            : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_io_hps_io_emac1_inst_RX_CTL                                         : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_hps_io_emac1_inst_TX_CTL                                         : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_io_hps_io_emac1_inst_RX_CLK                                         : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_hps_io_emac1_inst_RXD1                                           : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_hps_io_emac1_inst_RXD2                                           : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_hps_io_emac1_inst_RXD3                                           : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_hps_io_qspi_inst_IO0                                             : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO0
			hps_io_hps_io_qspi_inst_IO1                                             : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO1
			hps_io_hps_io_qspi_inst_IO2                                             : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO2
			hps_io_hps_io_qspi_inst_IO3                                             : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO3
			hps_io_hps_io_qspi_inst_SS0                                             : out   std_logic;                                        -- hps_io_qspi_inst_SS0
			hps_io_hps_io_qspi_inst_CLK                                             : out   std_logic;                                        -- hps_io_qspi_inst_CLK
			hps_io_hps_io_sdio_inst_CMD                                             : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_hps_io_sdio_inst_D0                                              : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_hps_io_sdio_inst_D1                                              : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_hps_io_sdio_inst_CLK                                             : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_hps_io_sdio_inst_D2                                              : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_hps_io_sdio_inst_D3                                              : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_hps_io_usb1_inst_D0                                              : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D0
			hps_io_hps_io_usb1_inst_D1                                              : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D1
			hps_io_hps_io_usb1_inst_D2                                              : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D2
			hps_io_hps_io_usb1_inst_D3                                              : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D3
			hps_io_hps_io_usb1_inst_D4                                              : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D4
			hps_io_hps_io_usb1_inst_D5                                              : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D5
			hps_io_hps_io_usb1_inst_D6                                              : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D6
			hps_io_hps_io_usb1_inst_D7                                              : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D7
			hps_io_hps_io_usb1_inst_CLK                                             : in    std_logic                     := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_hps_io_usb1_inst_STP                                             : out   std_logic;                                        -- hps_io_usb1_inst_STP
			hps_io_hps_io_usb1_inst_DIR                                             : in    std_logic                     := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_hps_io_usb1_inst_NXT                                             : in    std_logic                     := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_hps_io_spim1_inst_CLK                                            : out   std_logic;                                        -- hps_io_spim1_inst_CLK
			hps_io_hps_io_spim1_inst_MOSI                                           : out   std_logic;                                        -- hps_io_spim1_inst_MOSI
			hps_io_hps_io_spim1_inst_MISO                                           : in    std_logic                     := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_hps_io_spim1_inst_SS0                                            : out   std_logic;                                        -- hps_io_spim1_inst_SS0
			hps_io_hps_io_uart0_inst_RX                                             : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_hps_io_uart0_inst_TX                                             : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_io_hps_io_i2c0_inst_SDA                                             : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_hps_io_i2c0_inst_SCL                                             : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_hps_io_i2c1_inst_SDA                                             : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_hps_io_i2c1_inst_SCL                                             : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_hps_io_gpio_inst_GPIO09                                          : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_hps_io_gpio_inst_GPIO35                                          : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_hps_io_gpio_inst_GPIO40                                          : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_hps_io_gpio_inst_GPIO41                                          : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO41
			hps_io_hps_io_gpio_inst_GPIO48                                          : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO48
			hps_io_hps_io_gpio_inst_GPIO53                                          : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_hps_io_gpio_inst_GPIO54                                          : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_hps_io_gpio_inst_GPIO61                                          : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO61
			memory_mem_a                                                            : out   std_logic_vector(14 downto 0);                    -- mem_a
			memory_mem_ba                                                           : out   std_logic_vector(2 downto 0);                     -- mem_ba
			memory_mem_ck                                                           : out   std_logic;                                        -- mem_ck
			memory_mem_ck_n                                                         : out   std_logic;                                        -- mem_ck_n
			memory_mem_cke                                                          : out   std_logic;                                        -- mem_cke
			memory_mem_cs_n                                                         : out   std_logic;                                        -- mem_cs_n
			memory_mem_ras_n                                                        : out   std_logic;                                        -- mem_ras_n
			memory_mem_cas_n                                                        : out   std_logic;                                        -- mem_cas_n
			memory_mem_we_n                                                         : out   std_logic;                                        -- mem_we_n
			memory_mem_reset_n                                                      : out   std_logic;                                        -- mem_reset_n
			memory_mem_dq                                                           : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			memory_mem_dqs                                                          : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			memory_mem_dqs_n                                                        : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			memory_mem_odt                                                          : out   std_logic;                                        -- mem_odt
			memory_mem_dm                                                           : out   std_logic_vector(3 downto 0);                     -- mem_dm
			memory_oct_rzqin                                                        : in    std_logic                     := 'X';             -- oct_rzqin
			pixel_clk_clk                                                           : out   std_logic;                                        -- clk
			pll_vga_clk_25_clk                                                      : out   std_logic;                                        -- clk
			rgba_image_sink_data_valid                                              : in    std_logic                     := 'X';             -- data_valid
			rgba_image_sink_input_data                                              : in    std_logic_vector(31 downto 0) := (others => 'X'); -- input_data
			rgba_image_sink_img_width                                               : in    std_logic_vector(15 downto 0) := (others => 'X'); -- img_width
			rgba_image_sink_img_height                                              : in    std_logic_vector(15 downto 0) := (others => 'X'); -- img_height
			rgba_image_src_data                                                     : out   std_logic_vector(31 downto 0);                    -- data
			rgba_image_src_valid                                                    : out   std_logic;                                        -- valid
			rgba_stream_reset_reset_n                                               : in    std_logic                     := 'X';             -- reset_n
			sdram_ctrl_addr                                                         : out   std_logic_vector(12 downto 0);                    -- addr
			sdram_ctrl_ba                                                           : out   std_logic_vector(1 downto 0);                     -- ba
			sdram_ctrl_cas_n                                                        : out   std_logic;                                        -- cas_n
			sdram_ctrl_cke                                                          : out   std_logic;                                        -- cke
			sdram_ctrl_cs_n                                                         : out   std_logic;                                        -- cs_n
			sdram_ctrl_dq                                                           : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			sdram_ctrl_dqm                                                          : out   std_logic_vector(1 downto 0);                     -- dqm
			sdram_ctrl_ras_n                                                        : out   std_logic;                                        -- ras_n
			sdram_ctrl_we_n                                                         : out   std_logic;                                        -- we_n
			stream_control_endofpacket                                              : in    std_logic                     := 'X';             -- endofpacket
			stream_control_ready                                                    : out   std_logic;                                        -- ready
			stream_control_sreset                                                   : out   std_logic;                                        -- sreset
			stream_control_startofpacket                                            : in    std_logic                     := 'X';             -- startofpacket
			stream_control_frame_transition                                         : out   std_logic;                                        -- frame_transition
			system_pll_ref_clk_clk                                                  : in    std_logic                     := 'X';             -- clk
			system_pll_ref_reset_reset                                              : in    std_logic                     := 'X';             -- reset
			video_in_TD_CLK27                                                       : in    std_logic                     := 'X';             -- TD_CLK27
			video_in_TD_DATA                                                        : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- TD_DATA
			video_in_TD_HS                                                          : in    std_logic                     := 'X';             -- TD_HS
			video_in_TD_VS                                                          : in    std_logic                     := 'X';             -- TD_VS
			video_in_clk27_reset                                                    : in    std_logic                     := 'X';             -- clk27_reset
			video_in_TD_RESET                                                       : out   std_logic;                                        -- TD_RESET
			video_in_overflow_flag                                                  : out   std_logic;                                        -- overflow_flag
			video_subsystem_video_in_feed_forward_avalon_forward_sink_data          : in    std_logic_vector(23 downto 0) := (others => 'X'); -- data
			video_subsystem_video_in_feed_forward_avalon_forward_sink_startofpacket : in    std_logic                     := 'X';             -- startofpacket
			video_subsystem_video_in_feed_forward_avalon_forward_sink_endofpacket   : in    std_logic                     := 'X';             -- endofpacket
			video_subsystem_video_in_feed_forward_avalon_forward_sink_empty         : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			video_subsystem_video_in_feed_forward_avalon_forward_sink_valid         : in    std_logic                     := 'X';             -- valid
			video_subsystem_video_in_feed_forward_avalon_forward_sink_ready         : out   std_logic;                                        -- ready
			video_subsystem_video_in_scaler_avalon_scaler_source_ready              : in    std_logic                     := 'X';             -- ready
			video_subsystem_video_in_scaler_avalon_scaler_source_startofpacket      : out   std_logic;                                        -- startofpacket
			video_subsystem_video_in_scaler_avalon_scaler_source_endofpacket        : out   std_logic;                                        -- endofpacket
			video_subsystem_video_in_scaler_avalon_scaler_source_valid              : out   std_logic;                                        -- valid
			video_subsystem_video_in_scaler_avalon_scaler_source_data               : out   std_logic_vector(23 downto 0);                    -- data
			video_subsystem_video_in_scaler_avalon_scaler_source_channel            : out   std_logic                                         -- channel
		);
	end component Computer_System;

	u0 : component Computer_System
		port map (
			av_config_SDAT                                                          => CONNECTED_TO_av_config_SDAT,                                                          --                                                 av_config.SDAT
			av_config_SCLK                                                          => CONNECTED_TO_av_config_SCLK,                                                          --                                                          .SCLK
			h2f_reset_reset_n                                                       => CONNECTED_TO_h2f_reset_reset_n,                                                       --                                                 h2f_reset.reset_n
			hps_io_hps_io_emac1_inst_TX_CLK                                         => CONNECTED_TO_hps_io_hps_io_emac1_inst_TX_CLK,                                         --                                                    hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_hps_io_emac1_inst_TXD0                                           => CONNECTED_TO_hps_io_hps_io_emac1_inst_TXD0,                                           --                                                          .hps_io_emac1_inst_TXD0
			hps_io_hps_io_emac1_inst_TXD1                                           => CONNECTED_TO_hps_io_hps_io_emac1_inst_TXD1,                                           --                                                          .hps_io_emac1_inst_TXD1
			hps_io_hps_io_emac1_inst_TXD2                                           => CONNECTED_TO_hps_io_hps_io_emac1_inst_TXD2,                                           --                                                          .hps_io_emac1_inst_TXD2
			hps_io_hps_io_emac1_inst_TXD3                                           => CONNECTED_TO_hps_io_hps_io_emac1_inst_TXD3,                                           --                                                          .hps_io_emac1_inst_TXD3
			hps_io_hps_io_emac1_inst_RXD0                                           => CONNECTED_TO_hps_io_hps_io_emac1_inst_RXD0,                                           --                                                          .hps_io_emac1_inst_RXD0
			hps_io_hps_io_emac1_inst_MDIO                                           => CONNECTED_TO_hps_io_hps_io_emac1_inst_MDIO,                                           --                                                          .hps_io_emac1_inst_MDIO
			hps_io_hps_io_emac1_inst_MDC                                            => CONNECTED_TO_hps_io_hps_io_emac1_inst_MDC,                                            --                                                          .hps_io_emac1_inst_MDC
			hps_io_hps_io_emac1_inst_RX_CTL                                         => CONNECTED_TO_hps_io_hps_io_emac1_inst_RX_CTL,                                         --                                                          .hps_io_emac1_inst_RX_CTL
			hps_io_hps_io_emac1_inst_TX_CTL                                         => CONNECTED_TO_hps_io_hps_io_emac1_inst_TX_CTL,                                         --                                                          .hps_io_emac1_inst_TX_CTL
			hps_io_hps_io_emac1_inst_RX_CLK                                         => CONNECTED_TO_hps_io_hps_io_emac1_inst_RX_CLK,                                         --                                                          .hps_io_emac1_inst_RX_CLK
			hps_io_hps_io_emac1_inst_RXD1                                           => CONNECTED_TO_hps_io_hps_io_emac1_inst_RXD1,                                           --                                                          .hps_io_emac1_inst_RXD1
			hps_io_hps_io_emac1_inst_RXD2                                           => CONNECTED_TO_hps_io_hps_io_emac1_inst_RXD2,                                           --                                                          .hps_io_emac1_inst_RXD2
			hps_io_hps_io_emac1_inst_RXD3                                           => CONNECTED_TO_hps_io_hps_io_emac1_inst_RXD3,                                           --                                                          .hps_io_emac1_inst_RXD3
			hps_io_hps_io_qspi_inst_IO0                                             => CONNECTED_TO_hps_io_hps_io_qspi_inst_IO0,                                             --                                                          .hps_io_qspi_inst_IO0
			hps_io_hps_io_qspi_inst_IO1                                             => CONNECTED_TO_hps_io_hps_io_qspi_inst_IO1,                                             --                                                          .hps_io_qspi_inst_IO1
			hps_io_hps_io_qspi_inst_IO2                                             => CONNECTED_TO_hps_io_hps_io_qspi_inst_IO2,                                             --                                                          .hps_io_qspi_inst_IO2
			hps_io_hps_io_qspi_inst_IO3                                             => CONNECTED_TO_hps_io_hps_io_qspi_inst_IO3,                                             --                                                          .hps_io_qspi_inst_IO3
			hps_io_hps_io_qspi_inst_SS0                                             => CONNECTED_TO_hps_io_hps_io_qspi_inst_SS0,                                             --                                                          .hps_io_qspi_inst_SS0
			hps_io_hps_io_qspi_inst_CLK                                             => CONNECTED_TO_hps_io_hps_io_qspi_inst_CLK,                                             --                                                          .hps_io_qspi_inst_CLK
			hps_io_hps_io_sdio_inst_CMD                                             => CONNECTED_TO_hps_io_hps_io_sdio_inst_CMD,                                             --                                                          .hps_io_sdio_inst_CMD
			hps_io_hps_io_sdio_inst_D0                                              => CONNECTED_TO_hps_io_hps_io_sdio_inst_D0,                                              --                                                          .hps_io_sdio_inst_D0
			hps_io_hps_io_sdio_inst_D1                                              => CONNECTED_TO_hps_io_hps_io_sdio_inst_D1,                                              --                                                          .hps_io_sdio_inst_D1
			hps_io_hps_io_sdio_inst_CLK                                             => CONNECTED_TO_hps_io_hps_io_sdio_inst_CLK,                                             --                                                          .hps_io_sdio_inst_CLK
			hps_io_hps_io_sdio_inst_D2                                              => CONNECTED_TO_hps_io_hps_io_sdio_inst_D2,                                              --                                                          .hps_io_sdio_inst_D2
			hps_io_hps_io_sdio_inst_D3                                              => CONNECTED_TO_hps_io_hps_io_sdio_inst_D3,                                              --                                                          .hps_io_sdio_inst_D3
			hps_io_hps_io_usb1_inst_D0                                              => CONNECTED_TO_hps_io_hps_io_usb1_inst_D0,                                              --                                                          .hps_io_usb1_inst_D0
			hps_io_hps_io_usb1_inst_D1                                              => CONNECTED_TO_hps_io_hps_io_usb1_inst_D1,                                              --                                                          .hps_io_usb1_inst_D1
			hps_io_hps_io_usb1_inst_D2                                              => CONNECTED_TO_hps_io_hps_io_usb1_inst_D2,                                              --                                                          .hps_io_usb1_inst_D2
			hps_io_hps_io_usb1_inst_D3                                              => CONNECTED_TO_hps_io_hps_io_usb1_inst_D3,                                              --                                                          .hps_io_usb1_inst_D3
			hps_io_hps_io_usb1_inst_D4                                              => CONNECTED_TO_hps_io_hps_io_usb1_inst_D4,                                              --                                                          .hps_io_usb1_inst_D4
			hps_io_hps_io_usb1_inst_D5                                              => CONNECTED_TO_hps_io_hps_io_usb1_inst_D5,                                              --                                                          .hps_io_usb1_inst_D5
			hps_io_hps_io_usb1_inst_D6                                              => CONNECTED_TO_hps_io_hps_io_usb1_inst_D6,                                              --                                                          .hps_io_usb1_inst_D6
			hps_io_hps_io_usb1_inst_D7                                              => CONNECTED_TO_hps_io_hps_io_usb1_inst_D7,                                              --                                                          .hps_io_usb1_inst_D7
			hps_io_hps_io_usb1_inst_CLK                                             => CONNECTED_TO_hps_io_hps_io_usb1_inst_CLK,                                             --                                                          .hps_io_usb1_inst_CLK
			hps_io_hps_io_usb1_inst_STP                                             => CONNECTED_TO_hps_io_hps_io_usb1_inst_STP,                                             --                                                          .hps_io_usb1_inst_STP
			hps_io_hps_io_usb1_inst_DIR                                             => CONNECTED_TO_hps_io_hps_io_usb1_inst_DIR,                                             --                                                          .hps_io_usb1_inst_DIR
			hps_io_hps_io_usb1_inst_NXT                                             => CONNECTED_TO_hps_io_hps_io_usb1_inst_NXT,                                             --                                                          .hps_io_usb1_inst_NXT
			hps_io_hps_io_spim1_inst_CLK                                            => CONNECTED_TO_hps_io_hps_io_spim1_inst_CLK,                                            --                                                          .hps_io_spim1_inst_CLK
			hps_io_hps_io_spim1_inst_MOSI                                           => CONNECTED_TO_hps_io_hps_io_spim1_inst_MOSI,                                           --                                                          .hps_io_spim1_inst_MOSI
			hps_io_hps_io_spim1_inst_MISO                                           => CONNECTED_TO_hps_io_hps_io_spim1_inst_MISO,                                           --                                                          .hps_io_spim1_inst_MISO
			hps_io_hps_io_spim1_inst_SS0                                            => CONNECTED_TO_hps_io_hps_io_spim1_inst_SS0,                                            --                                                          .hps_io_spim1_inst_SS0
			hps_io_hps_io_uart0_inst_RX                                             => CONNECTED_TO_hps_io_hps_io_uart0_inst_RX,                                             --                                                          .hps_io_uart0_inst_RX
			hps_io_hps_io_uart0_inst_TX                                             => CONNECTED_TO_hps_io_hps_io_uart0_inst_TX,                                             --                                                          .hps_io_uart0_inst_TX
			hps_io_hps_io_i2c0_inst_SDA                                             => CONNECTED_TO_hps_io_hps_io_i2c0_inst_SDA,                                             --                                                          .hps_io_i2c0_inst_SDA
			hps_io_hps_io_i2c0_inst_SCL                                             => CONNECTED_TO_hps_io_hps_io_i2c0_inst_SCL,                                             --                                                          .hps_io_i2c0_inst_SCL
			hps_io_hps_io_i2c1_inst_SDA                                             => CONNECTED_TO_hps_io_hps_io_i2c1_inst_SDA,                                             --                                                          .hps_io_i2c1_inst_SDA
			hps_io_hps_io_i2c1_inst_SCL                                             => CONNECTED_TO_hps_io_hps_io_i2c1_inst_SCL,                                             --                                                          .hps_io_i2c1_inst_SCL
			hps_io_hps_io_gpio_inst_GPIO09                                          => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO09,                                          --                                                          .hps_io_gpio_inst_GPIO09
			hps_io_hps_io_gpio_inst_GPIO35                                          => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO35,                                          --                                                          .hps_io_gpio_inst_GPIO35
			hps_io_hps_io_gpio_inst_GPIO40                                          => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO40,                                          --                                                          .hps_io_gpio_inst_GPIO40
			hps_io_hps_io_gpio_inst_GPIO41                                          => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO41,                                          --                                                          .hps_io_gpio_inst_GPIO41
			hps_io_hps_io_gpio_inst_GPIO48                                          => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO48,                                          --                                                          .hps_io_gpio_inst_GPIO48
			hps_io_hps_io_gpio_inst_GPIO53                                          => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO53,                                          --                                                          .hps_io_gpio_inst_GPIO53
			hps_io_hps_io_gpio_inst_GPIO54                                          => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO54,                                          --                                                          .hps_io_gpio_inst_GPIO54
			hps_io_hps_io_gpio_inst_GPIO61                                          => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO61,                                          --                                                          .hps_io_gpio_inst_GPIO61
			memory_mem_a                                                            => CONNECTED_TO_memory_mem_a,                                                            --                                                    memory.mem_a
			memory_mem_ba                                                           => CONNECTED_TO_memory_mem_ba,                                                           --                                                          .mem_ba
			memory_mem_ck                                                           => CONNECTED_TO_memory_mem_ck,                                                           --                                                          .mem_ck
			memory_mem_ck_n                                                         => CONNECTED_TO_memory_mem_ck_n,                                                         --                                                          .mem_ck_n
			memory_mem_cke                                                          => CONNECTED_TO_memory_mem_cke,                                                          --                                                          .mem_cke
			memory_mem_cs_n                                                         => CONNECTED_TO_memory_mem_cs_n,                                                         --                                                          .mem_cs_n
			memory_mem_ras_n                                                        => CONNECTED_TO_memory_mem_ras_n,                                                        --                                                          .mem_ras_n
			memory_mem_cas_n                                                        => CONNECTED_TO_memory_mem_cas_n,                                                        --                                                          .mem_cas_n
			memory_mem_we_n                                                         => CONNECTED_TO_memory_mem_we_n,                                                         --                                                          .mem_we_n
			memory_mem_reset_n                                                      => CONNECTED_TO_memory_mem_reset_n,                                                      --                                                          .mem_reset_n
			memory_mem_dq                                                           => CONNECTED_TO_memory_mem_dq,                                                           --                                                          .mem_dq
			memory_mem_dqs                                                          => CONNECTED_TO_memory_mem_dqs,                                                          --                                                          .mem_dqs
			memory_mem_dqs_n                                                        => CONNECTED_TO_memory_mem_dqs_n,                                                        --                                                          .mem_dqs_n
			memory_mem_odt                                                          => CONNECTED_TO_memory_mem_odt,                                                          --                                                          .mem_odt
			memory_mem_dm                                                           => CONNECTED_TO_memory_mem_dm,                                                           --                                                          .mem_dm
			memory_oct_rzqin                                                        => CONNECTED_TO_memory_oct_rzqin,                                                        --                                                          .oct_rzqin
			pixel_clk_clk                                                           => CONNECTED_TO_pixel_clk_clk,                                                           --                                                 pixel_clk.clk
			pll_vga_clk_25_clk                                                      => CONNECTED_TO_pll_vga_clk_25_clk,                                                      --                                            pll_vga_clk_25.clk
			rgba_image_sink_data_valid                                              => CONNECTED_TO_rgba_image_sink_data_valid,                                              --                                           rgba_image_sink.data_valid
			rgba_image_sink_input_data                                              => CONNECTED_TO_rgba_image_sink_input_data,                                              --                                                          .input_data
			rgba_image_sink_img_width                                               => CONNECTED_TO_rgba_image_sink_img_width,                                               --                                                          .img_width
			rgba_image_sink_img_height                                              => CONNECTED_TO_rgba_image_sink_img_height,                                              --                                                          .img_height
			rgba_image_src_data                                                     => CONNECTED_TO_rgba_image_src_data,                                                     --                                            rgba_image_src.data
			rgba_image_src_valid                                                    => CONNECTED_TO_rgba_image_src_valid,                                                    --                                                          .valid
			rgba_stream_reset_reset_n                                               => CONNECTED_TO_rgba_stream_reset_reset_n,                                               --                                         rgba_stream_reset.reset_n
			sdram_ctrl_addr                                                         => CONNECTED_TO_sdram_ctrl_addr,                                                         --                                                sdram_ctrl.addr
			sdram_ctrl_ba                                                           => CONNECTED_TO_sdram_ctrl_ba,                                                           --                                                          .ba
			sdram_ctrl_cas_n                                                        => CONNECTED_TO_sdram_ctrl_cas_n,                                                        --                                                          .cas_n
			sdram_ctrl_cke                                                          => CONNECTED_TO_sdram_ctrl_cke,                                                          --                                                          .cke
			sdram_ctrl_cs_n                                                         => CONNECTED_TO_sdram_ctrl_cs_n,                                                         --                                                          .cs_n
			sdram_ctrl_dq                                                           => CONNECTED_TO_sdram_ctrl_dq,                                                           --                                                          .dq
			sdram_ctrl_dqm                                                          => CONNECTED_TO_sdram_ctrl_dqm,                                                          --                                                          .dqm
			sdram_ctrl_ras_n                                                        => CONNECTED_TO_sdram_ctrl_ras_n,                                                        --                                                          .ras_n
			sdram_ctrl_we_n                                                         => CONNECTED_TO_sdram_ctrl_we_n,                                                         --                                                          .we_n
			stream_control_endofpacket                                              => CONNECTED_TO_stream_control_endofpacket,                                              --                                            stream_control.endofpacket
			stream_control_ready                                                    => CONNECTED_TO_stream_control_ready,                                                    --                                                          .ready
			stream_control_sreset                                                   => CONNECTED_TO_stream_control_sreset,                                                   --                                                          .sreset
			stream_control_startofpacket                                            => CONNECTED_TO_stream_control_startofpacket,                                            --                                                          .startofpacket
			stream_control_frame_transition                                         => CONNECTED_TO_stream_control_frame_transition,                                         --                                                          .frame_transition
			system_pll_ref_clk_clk                                                  => CONNECTED_TO_system_pll_ref_clk_clk,                                                  --                                        system_pll_ref_clk.clk
			system_pll_ref_reset_reset                                              => CONNECTED_TO_system_pll_ref_reset_reset,                                              --                                      system_pll_ref_reset.reset
			video_in_TD_CLK27                                                       => CONNECTED_TO_video_in_TD_CLK27,                                                       --                                                  video_in.TD_CLK27
			video_in_TD_DATA                                                        => CONNECTED_TO_video_in_TD_DATA,                                                        --                                                          .TD_DATA
			video_in_TD_HS                                                          => CONNECTED_TO_video_in_TD_HS,                                                          --                                                          .TD_HS
			video_in_TD_VS                                                          => CONNECTED_TO_video_in_TD_VS,                                                          --                                                          .TD_VS
			video_in_clk27_reset                                                    => CONNECTED_TO_video_in_clk27_reset,                                                    --                                                          .clk27_reset
			video_in_TD_RESET                                                       => CONNECTED_TO_video_in_TD_RESET,                                                       --                                                          .TD_RESET
			video_in_overflow_flag                                                  => CONNECTED_TO_video_in_overflow_flag,                                                  --                                                          .overflow_flag
			video_subsystem_video_in_feed_forward_avalon_forward_sink_data          => CONNECTED_TO_video_subsystem_video_in_feed_forward_avalon_forward_sink_data,          -- video_subsystem_video_in_feed_forward_avalon_forward_sink.data
			video_subsystem_video_in_feed_forward_avalon_forward_sink_startofpacket => CONNECTED_TO_video_subsystem_video_in_feed_forward_avalon_forward_sink_startofpacket, --                                                          .startofpacket
			video_subsystem_video_in_feed_forward_avalon_forward_sink_endofpacket   => CONNECTED_TO_video_subsystem_video_in_feed_forward_avalon_forward_sink_endofpacket,   --                                                          .endofpacket
			video_subsystem_video_in_feed_forward_avalon_forward_sink_empty         => CONNECTED_TO_video_subsystem_video_in_feed_forward_avalon_forward_sink_empty,         --                                                          .empty
			video_subsystem_video_in_feed_forward_avalon_forward_sink_valid         => CONNECTED_TO_video_subsystem_video_in_feed_forward_avalon_forward_sink_valid,         --                                                          .valid
			video_subsystem_video_in_feed_forward_avalon_forward_sink_ready         => CONNECTED_TO_video_subsystem_video_in_feed_forward_avalon_forward_sink_ready,         --                                                          .ready
			video_subsystem_video_in_scaler_avalon_scaler_source_ready              => CONNECTED_TO_video_subsystem_video_in_scaler_avalon_scaler_source_ready,              --      video_subsystem_video_in_scaler_avalon_scaler_source.ready
			video_subsystem_video_in_scaler_avalon_scaler_source_startofpacket      => CONNECTED_TO_video_subsystem_video_in_scaler_avalon_scaler_source_startofpacket,      --                                                          .startofpacket
			video_subsystem_video_in_scaler_avalon_scaler_source_endofpacket        => CONNECTED_TO_video_subsystem_video_in_scaler_avalon_scaler_source_endofpacket,        --                                                          .endofpacket
			video_subsystem_video_in_scaler_avalon_scaler_source_valid              => CONNECTED_TO_video_subsystem_video_in_scaler_avalon_scaler_source_valid,              --                                                          .valid
			video_subsystem_video_in_scaler_avalon_scaler_source_data               => CONNECTED_TO_video_subsystem_video_in_scaler_avalon_scaler_source_data,               --                                                          .data
			video_subsystem_video_in_scaler_avalon_scaler_source_channel            => CONNECTED_TO_video_subsystem_video_in_scaler_avalon_scaler_source_channel             --                                                          .channel
		);

